/*********************************************/
/* SINE table of size 4096 and 13-bit values */
/* Latency: 4 CLK cycles                     */
/* TESTBENCH                                 */
/*********************************************/
`timescale 1ns / 1ps
module sin_cos_table_4096_13bit_tb ();

localparam     DATA_WIDTH = 13;
localparam     ADDR_WIDTH = 12;


    logic [15:0] cycleCounter = 0;
    logic CLK;
    logic CE;
    logic RESET;
    logic [ADDR_WIDTH-1:0] PHASE;
    wire signed [DATA_WIDTH-1:0] SIN_VALUE;
    wire signed [DATA_WIDTH-1:0] COS_VALUE;
    
    sin_cos_table_4096_13bit
    #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH)
    )
    sin_table_instance
    (
        .*
    );
    
    // drive CLK
    always begin
        #1.472 CLK=0;
        #1.472 CLK=1; 
        cycleCounter = cycleCounter + 1;
    end
    
    task nextCycle(input [ADDR_WIDTH-1:0] phase);
         begin
             @(posedge CLK) #1 ;
             PHASE = phase;
             $display("    [%d]   nextCycle PHASE=%d", cycleCounter, PHASE);
         end
    endtask
     
    task checkResult(input signed [DATA_WIDTH-1:0] expected_sin_value, input signed [DATA_WIDTH-1:0] expected_cos_value);
         begin
             $display("    [%d]             SIN=%d COS=%d", cycleCounter, SIN_VALUE, COS_VALUE);
             if (SIN_VALUE != expected_sin_value) begin
                 $display("    [%d] ERROR: SIN_VALUE does not match with expected result, expected %x actual %x", cycleCounter, expected_sin_value, SIN_VALUE);
                 $finish();
             end
             if (COS_VALUE != expected_cos_value) begin
                 $display("    [%d] ERROR: COS_VALUE does not match with expected result, expected %x actual %x", cycleCounter, expected_cos_value, COS_VALUE);
                 $finish();
             end
         end
    endtask
     
    // reset condition
    initial begin
        RESET = 0;
        CE = 0;
        #200 @(posedge CLK) RESET = 1;
        #100 @(posedge CLK) RESET = 0;
        @(posedge CLK) #1 CE = 1;
        PHASE = 0;
     
        $display("Starting verification");
    

        /* Outputs are delayed by 4 clock cycles */
        nextCycle(0);
        nextCycle(1);
        nextCycle(2);
        nextCycle(3);
        nextCycle(4); checkResult(3, 4095);
        nextCycle(5); checkResult(9, 4095);
        nextCycle(6); checkResult(16, 4095);
        nextCycle(7); checkResult(22, 4095);
        nextCycle(8); checkResult(28, 4095);
        nextCycle(9); checkResult(35, 4095);
        nextCycle(10); checkResult(41, 4095);
        nextCycle(11); checkResult(47, 4095);
        nextCycle(12); checkResult(53, 4095);
        nextCycle(13); checkResult(60, 4095);
        nextCycle(14); checkResult(66, 4094);
        nextCycle(15); checkResult(72, 4094);
        nextCycle(16); checkResult(79, 4094);
        nextCycle(17); checkResult(85, 4094);
        nextCycle(18); checkResult(91, 4094);
        nextCycle(19); checkResult(97, 4094);
        nextCycle(20); checkResult(104, 4094);
        nextCycle(21); checkResult(110, 4094);
        nextCycle(22); checkResult(116, 4093);
        nextCycle(23); checkResult(122, 4093);
        nextCycle(24); checkResult(129, 4093);
        nextCycle(25); checkResult(135, 4093);
        nextCycle(26); checkResult(141, 4093);
        nextCycle(27); checkResult(148, 4092);
        nextCycle(28); checkResult(154, 4092);
        nextCycle(29); checkResult(160, 4092);
        nextCycle(30); checkResult(166, 4092);
        nextCycle(31); checkResult(173, 4091);
        nextCycle(32); checkResult(179, 4091);
        nextCycle(33); checkResult(185, 4091);
        nextCycle(34); checkResult(192, 4091);
        nextCycle(35); checkResult(198, 4090);
        nextCycle(36); checkResult(204, 4090);
        nextCycle(37); checkResult(210, 4090);
        nextCycle(38); checkResult(217, 4089);
        nextCycle(39); checkResult(223, 4089);
        nextCycle(40); checkResult(229, 4089);
        nextCycle(41); checkResult(235, 4088);
        nextCycle(42); checkResult(242, 4088);
        nextCycle(43); checkResult(248, 4087);
        nextCycle(44); checkResult(254, 4087);
        nextCycle(45); checkResult(261, 4087);
        nextCycle(46); checkResult(267, 4086);
        nextCycle(47); checkResult(273, 4086);
        nextCycle(48); checkResult(279, 4085);
        nextCycle(49); checkResult(286, 4085);
        nextCycle(50); checkResult(292, 4085);
        nextCycle(51); checkResult(298, 4084);
        nextCycle(52); checkResult(304, 4084);
        nextCycle(53); checkResult(311, 4083);
        nextCycle(54); checkResult(317, 4083);
        nextCycle(55); checkResult(323, 4082);
        nextCycle(56); checkResult(329, 4082);
        nextCycle(57); checkResult(336, 4081);
        nextCycle(58); checkResult(342, 4081);
        nextCycle(59); checkResult(348, 4080);
        nextCycle(60); checkResult(354, 4080);
        nextCycle(61); checkResult(361, 4079);
        nextCycle(62); checkResult(367, 4079);
        nextCycle(63); checkResult(373, 4078);
        nextCycle(64); checkResult(379, 4077);
        nextCycle(65); checkResult(386, 4077);
        nextCycle(66); checkResult(392, 4076);
        nextCycle(67); checkResult(398, 4076);
        nextCycle(68); checkResult(405, 4075);
        nextCycle(69); checkResult(411, 4074);
        nextCycle(70); checkResult(417, 4074);
        nextCycle(71); checkResult(423, 4073);
        nextCycle(72); checkResult(430, 4072);
        nextCycle(73); checkResult(436, 4072);
        nextCycle(74); checkResult(442, 4071);
        nextCycle(75); checkResult(448, 4070);
        nextCycle(76); checkResult(454, 4070);
        nextCycle(77); checkResult(461, 4069);
        nextCycle(78); checkResult(467, 4068);
        nextCycle(79); checkResult(473, 4068);
        nextCycle(80); checkResult(479, 4067);
        nextCycle(81); checkResult(486, 4066);
        nextCycle(82); checkResult(492, 4065);
        nextCycle(83); checkResult(498, 4065);
        nextCycle(84); checkResult(504, 4064);
        nextCycle(85); checkResult(511, 4063);
        nextCycle(86); checkResult(517, 4062);
        nextCycle(87); checkResult(523, 4061);
        nextCycle(88); checkResult(529, 4061);
        nextCycle(89); checkResult(536, 4060);
        nextCycle(90); checkResult(542, 4059);
        nextCycle(91); checkResult(548, 4058);
        nextCycle(92); checkResult(554, 4057);
        nextCycle(93); checkResult(560, 4056);
        nextCycle(94); checkResult(567, 4056);
        nextCycle(95); checkResult(573, 4055);
        nextCycle(96); checkResult(579, 4054);
        nextCycle(97); checkResult(585, 4053);
        nextCycle(98); checkResult(592, 4052);
        nextCycle(99); checkResult(598, 4051);
        nextCycle(100); checkResult(604, 4050);
        nextCycle(101); checkResult(610, 4049);
        nextCycle(102); checkResult(616, 4048);
        nextCycle(103); checkResult(623, 4047);
        nextCycle(104); checkResult(629, 4046);
        nextCycle(105); checkResult(635, 4045);
        nextCycle(106); checkResult(641, 4044);
        nextCycle(107); checkResult(647, 4043);
        nextCycle(108); checkResult(654, 4042);
        nextCycle(109); checkResult(660, 4041);
        nextCycle(110); checkResult(666, 4040);
        nextCycle(111); checkResult(672, 4039);
        nextCycle(112); checkResult(678, 4038);
        nextCycle(113); checkResult(685, 4037);
        nextCycle(114); checkResult(691, 4036);
        nextCycle(115); checkResult(697, 4035);
        nextCycle(116); checkResult(703, 4034);
        nextCycle(117); checkResult(709, 4033);
        nextCycle(118); checkResult(716, 4032);
        nextCycle(119); checkResult(722, 4031);
        nextCycle(120); checkResult(728, 4030);
        nextCycle(121); checkResult(734, 4029);
        nextCycle(122); checkResult(740, 4028);
        nextCycle(123); checkResult(746, 4026);
        nextCycle(124); checkResult(753, 4025);
        nextCycle(125); checkResult(759, 4024);
        nextCycle(126); checkResult(765, 4023);
        nextCycle(127); checkResult(771, 4022);
        nextCycle(128); checkResult(777, 4021);
        nextCycle(129); checkResult(783, 4019);
        nextCycle(130); checkResult(790, 4018);
        nextCycle(131); checkResult(796, 4017);
        nextCycle(132); checkResult(802, 4016);
        nextCycle(133); checkResult(808, 4014);
        nextCycle(134); checkResult(814, 4013);
        nextCycle(135); checkResult(820, 4012);
        nextCycle(136); checkResult(827, 4011);
        nextCycle(137); checkResult(833, 4009);
        nextCycle(138); checkResult(839, 4008);
        nextCycle(139); checkResult(845, 4007);
        nextCycle(140); checkResult(851, 4006);
        nextCycle(141); checkResult(857, 4004);
        nextCycle(142); checkResult(863, 4003);
        nextCycle(143); checkResult(870, 4002);
        nextCycle(144); checkResult(876, 4000);
        nextCycle(145); checkResult(882, 3999);
        nextCycle(146); checkResult(888, 3998);
        nextCycle(147); checkResult(894, 3996);
        nextCycle(148); checkResult(900, 3995);
        nextCycle(149); checkResult(906, 3993);
        nextCycle(150); checkResult(913, 3992);
        nextCycle(151); checkResult(919, 3991);
        nextCycle(152); checkResult(925, 3989);
        nextCycle(153); checkResult(931, 3988);
        nextCycle(154); checkResult(937, 3986);
        nextCycle(155); checkResult(943, 3985);
        nextCycle(156); checkResult(949, 3983);
        nextCycle(157); checkResult(955, 3982);
        nextCycle(158); checkResult(961, 3981);
        nextCycle(159); checkResult(968, 3979);
        nextCycle(160); checkResult(974, 3978);
        nextCycle(161); checkResult(980, 3976);
        nextCycle(162); checkResult(986, 3975);
        nextCycle(163); checkResult(992, 3973);
        nextCycle(164); checkResult(998, 3972);
        nextCycle(165); checkResult(1004, 3970);
        nextCycle(166); checkResult(1010, 3968);
        nextCycle(167); checkResult(1016, 3967);
        nextCycle(168); checkResult(1022, 3965);
        nextCycle(169); checkResult(1028, 3964);
        nextCycle(170); checkResult(1035, 3962);
        nextCycle(171); checkResult(1041, 3961);
        nextCycle(172); checkResult(1047, 3959);
        nextCycle(173); checkResult(1053, 3957);
        nextCycle(174); checkResult(1059, 3956);
        nextCycle(175); checkResult(1065, 3954);
        nextCycle(176); checkResult(1071, 3952);
        nextCycle(177); checkResult(1077, 3951);
        nextCycle(178); checkResult(1083, 3949);
        nextCycle(179); checkResult(1089, 3947);
        nextCycle(180); checkResult(1095, 3946);
        nextCycle(181); checkResult(1101, 3944);
        nextCycle(182); checkResult(1107, 3942);
        nextCycle(183); checkResult(1113, 3941);
        nextCycle(184); checkResult(1119, 3939);
        nextCycle(185); checkResult(1125, 3937);
        nextCycle(186); checkResult(1131, 3936);
        nextCycle(187); checkResult(1138, 3934);
        nextCycle(188); checkResult(1144, 3932);
        nextCycle(189); checkResult(1150, 3930);
        nextCycle(190); checkResult(1156, 3929);
        nextCycle(191); checkResult(1162, 3927);
        nextCycle(192); checkResult(1168, 3925);
        nextCycle(193); checkResult(1174, 3923);
        nextCycle(194); checkResult(1180, 3921);
        nextCycle(195); checkResult(1186, 3920);
        nextCycle(196); checkResult(1192, 3918);
        nextCycle(197); checkResult(1198, 3916);
        nextCycle(198); checkResult(1204, 3914);
        nextCycle(199); checkResult(1210, 3912);
        nextCycle(200); checkResult(1216, 3910);
        nextCycle(201); checkResult(1222, 3909);
        nextCycle(202); checkResult(1228, 3907);
        nextCycle(203); checkResult(1234, 3905);
        nextCycle(204); checkResult(1240, 3903);
        nextCycle(205); checkResult(1246, 3901);
        nextCycle(206); checkResult(1252, 3899);
        nextCycle(207); checkResult(1258, 3897);
        nextCycle(208); checkResult(1264, 3895);
        nextCycle(209); checkResult(1270, 3893);
        nextCycle(210); checkResult(1276, 3891);
        nextCycle(211); checkResult(1282, 3889);
        nextCycle(212); checkResult(1288, 3887);
        nextCycle(213); checkResult(1293, 3885);
        nextCycle(214); checkResult(1299, 3883);
        nextCycle(215); checkResult(1305, 3881);
        nextCycle(216); checkResult(1311, 3879);
        nextCycle(217); checkResult(1317, 3877);
        nextCycle(218); checkResult(1323, 3875);
        nextCycle(219); checkResult(1329, 3873);
        nextCycle(220); checkResult(1335, 3871);
        nextCycle(221); checkResult(1341, 3869);
        nextCycle(222); checkResult(1347, 3867);
        nextCycle(223); checkResult(1353, 3865);
        nextCycle(224); checkResult(1359, 3863);
        nextCycle(225); checkResult(1365, 3861);
        nextCycle(226); checkResult(1371, 3859);
        nextCycle(227); checkResult(1377, 3857);
        nextCycle(228); checkResult(1383, 3855);
        nextCycle(229); checkResult(1388, 3852);
        nextCycle(230); checkResult(1394, 3850);
        nextCycle(231); checkResult(1400, 3848);
        nextCycle(232); checkResult(1406, 3846);
        nextCycle(233); checkResult(1412, 3844);
        nextCycle(234); checkResult(1418, 3842);
        nextCycle(235); checkResult(1424, 3839);
        nextCycle(236); checkResult(1430, 3837);
        nextCycle(237); checkResult(1436, 3835);
        nextCycle(238); checkResult(1441, 3833);
        nextCycle(239); checkResult(1447, 3831);
        nextCycle(240); checkResult(1453, 3828);
        nextCycle(241); checkResult(1459, 3826);
        nextCycle(242); checkResult(1465, 3824);
        nextCycle(243); checkResult(1471, 3822);
        nextCycle(244); checkResult(1477, 3819);
        nextCycle(245); checkResult(1483, 3817);
        nextCycle(246); checkResult(1488, 3815);
        nextCycle(247); checkResult(1494, 3813);
        nextCycle(248); checkResult(1500, 3810);
        nextCycle(249); checkResult(1506, 3808);
        nextCycle(250); checkResult(1512, 3806);
        nextCycle(251); checkResult(1518, 3803);
        nextCycle(252); checkResult(1523, 3801);
        nextCycle(253); checkResult(1529, 3799);
        nextCycle(254); checkResult(1535, 3796);
        nextCycle(255); checkResult(1541, 3794);
        nextCycle(256); checkResult(1547, 3792);
        nextCycle(257); checkResult(1553, 3789);
        nextCycle(258); checkResult(1558, 3787);
        nextCycle(259); checkResult(1564, 3784);
        nextCycle(260); checkResult(1570, 3782);
        nextCycle(261); checkResult(1576, 3780);
        nextCycle(262); checkResult(1582, 3777);
        nextCycle(263); checkResult(1587, 3775);
        nextCycle(264); checkResult(1593, 3772);
        nextCycle(265); checkResult(1599, 3770);
        nextCycle(266); checkResult(1605, 3767);
        nextCycle(267); checkResult(1611, 3765);
        nextCycle(268); checkResult(1616, 3763);
        nextCycle(269); checkResult(1622, 3760);
        nextCycle(270); checkResult(1628, 3758);
        nextCycle(271); checkResult(1634, 3755);
        nextCycle(272); checkResult(1639, 3753);
        nextCycle(273); checkResult(1645, 3750);
        nextCycle(274); checkResult(1651, 3747);
        nextCycle(275); checkResult(1657, 3745);
        nextCycle(276); checkResult(1662, 3742);
        nextCycle(277); checkResult(1668, 3740);
        nextCycle(278); checkResult(1674, 3737);
        nextCycle(279); checkResult(1680, 3735);
        nextCycle(280); checkResult(1685, 3732);
        nextCycle(281); checkResult(1691, 3730);
        nextCycle(282); checkResult(1697, 3727);
        nextCycle(283); checkResult(1702, 3724);
        nextCycle(284); checkResult(1708, 3722);
        nextCycle(285); checkResult(1714, 3719);
        nextCycle(286); checkResult(1720, 3716);
        nextCycle(287); checkResult(1725, 3714);
        nextCycle(288); checkResult(1731, 3711);
        nextCycle(289); checkResult(1737, 3709);
        nextCycle(290); checkResult(1742, 3706);
        nextCycle(291); checkResult(1748, 3703);
        nextCycle(292); checkResult(1754, 3700);
        nextCycle(293); checkResult(1759, 3698);
        nextCycle(294); checkResult(1765, 3695);
        nextCycle(295); checkResult(1771, 3692);
        nextCycle(296); checkResult(1776, 3690);
        nextCycle(297); checkResult(1782, 3687);
        nextCycle(298); checkResult(1788, 3684);
        nextCycle(299); checkResult(1793, 3681);
        nextCycle(300); checkResult(1799, 3679);
        nextCycle(301); checkResult(1805, 3676);
        nextCycle(302); checkResult(1810, 3673);
        nextCycle(303); checkResult(1816, 3670);
        nextCycle(304); checkResult(1821, 3668);
        nextCycle(305); checkResult(1827, 3665);
        nextCycle(306); checkResult(1833, 3662);
        nextCycle(307); checkResult(1838, 3659);
        nextCycle(308); checkResult(1844, 3656);
        nextCycle(309); checkResult(1850, 3654);
        nextCycle(310); checkResult(1855, 3651);
        nextCycle(311); checkResult(1861, 3648);
        nextCycle(312); checkResult(1866, 3645);
        nextCycle(313); checkResult(1872, 3642);
        nextCycle(314); checkResult(1878, 3639);
        nextCycle(315); checkResult(1883, 3636);
        nextCycle(316); checkResult(1889, 3633);
        nextCycle(317); checkResult(1894, 3631);
        nextCycle(318); checkResult(1900, 3628);
        nextCycle(319); checkResult(1905, 3625);
        nextCycle(320); checkResult(1911, 3622);
        nextCycle(321); checkResult(1917, 3619);
        nextCycle(322); checkResult(1922, 3616);
        nextCycle(323); checkResult(1928, 3613);
        nextCycle(324); checkResult(1933, 3610);
        nextCycle(325); checkResult(1939, 3607);
        nextCycle(326); checkResult(1944, 3604);
        nextCycle(327); checkResult(1950, 3601);
        nextCycle(328); checkResult(1955, 3598);
        nextCycle(329); checkResult(1961, 3595);
        nextCycle(330); checkResult(1966, 3592);
        nextCycle(331); checkResult(1972, 3589);
        nextCycle(332); checkResult(1977, 3586);
        nextCycle(333); checkResult(1983, 3583);
        nextCycle(334); checkResult(1988, 3580);
        nextCycle(335); checkResult(1994, 3577);
        nextCycle(336); checkResult(1999, 3574);
        nextCycle(337); checkResult(2005, 3571);
        nextCycle(338); checkResult(2010, 3568);
        nextCycle(339); checkResult(2016, 3565);
        nextCycle(340); checkResult(2021, 3561);
        nextCycle(341); checkResult(2027, 3558);
        nextCycle(342); checkResult(2032, 3555);
        nextCycle(343); checkResult(2038, 3552);
        nextCycle(344); checkResult(2043, 3549);
        nextCycle(345); checkResult(2048, 3546);
        nextCycle(346); checkResult(2054, 3543);
        nextCycle(347); checkResult(2059, 3540);
        nextCycle(348); checkResult(2065, 3536);
        nextCycle(349); checkResult(2070, 3533);
        nextCycle(350); checkResult(2076, 3530);
        nextCycle(351); checkResult(2081, 3527);
        nextCycle(352); checkResult(2086, 3524);
        nextCycle(353); checkResult(2092, 3520);
        nextCycle(354); checkResult(2097, 3517);
        nextCycle(355); checkResult(2103, 3514);
        nextCycle(356); checkResult(2108, 3511);
        nextCycle(357); checkResult(2113, 3508);
        nextCycle(358); checkResult(2119, 3504);
        nextCycle(359); checkResult(2124, 3501);
        nextCycle(360); checkResult(2129, 3498);
        nextCycle(361); checkResult(2135, 3495);
        nextCycle(362); checkResult(2140, 3491);
        nextCycle(363); checkResult(2146, 3488);
        nextCycle(364); checkResult(2151, 3485);
        nextCycle(365); checkResult(2156, 3481);
        nextCycle(366); checkResult(2162, 3478);
        nextCycle(367); checkResult(2167, 3475);
        nextCycle(368); checkResult(2172, 3471);
        nextCycle(369); checkResult(2178, 3468);
        nextCycle(370); checkResult(2183, 3465);
        nextCycle(371); checkResult(2188, 3461);
        nextCycle(372); checkResult(2193, 3458);
        nextCycle(373); checkResult(2199, 3455);
        nextCycle(374); checkResult(2204, 3451);
        nextCycle(375); checkResult(2209, 3448);
        nextCycle(376); checkResult(2215, 3444);
        nextCycle(377); checkResult(2220, 3441);
        nextCycle(378); checkResult(2225, 3438);
        nextCycle(379); checkResult(2230, 3434);
        nextCycle(380); checkResult(2236, 3431);
        nextCycle(381); checkResult(2241, 3427);
        nextCycle(382); checkResult(2246, 3424);
        nextCycle(383); checkResult(2252, 3420);
        nextCycle(384); checkResult(2257, 3417);
        nextCycle(385); checkResult(2262, 3414);
        nextCycle(386); checkResult(2267, 3410);
        nextCycle(387); checkResult(2272, 3407);
        nextCycle(388); checkResult(2278, 3403);
        nextCycle(389); checkResult(2283, 3400);
        nextCycle(390); checkResult(2288, 3396);
        nextCycle(391); checkResult(2293, 3393);
        nextCycle(392); checkResult(2299, 3389);
        nextCycle(393); checkResult(2304, 3386);
        nextCycle(394); checkResult(2309, 3382);
        nextCycle(395); checkResult(2314, 3378);
        nextCycle(396); checkResult(2319, 3375);
        nextCycle(397); checkResult(2324, 3371);
        nextCycle(398); checkResult(2330, 3368);
        nextCycle(399); checkResult(2335, 3364);
        nextCycle(400); checkResult(2340, 3361);
        nextCycle(401); checkResult(2345, 3357);
        nextCycle(402); checkResult(2350, 3353);
        nextCycle(403); checkResult(2355, 3350);
        nextCycle(404); checkResult(2361, 3346);
        nextCycle(405); checkResult(2366, 3343);
        nextCycle(406); checkResult(2371, 3339);
        nextCycle(407); checkResult(2376, 3335);
        nextCycle(408); checkResult(2381, 3332);
        nextCycle(409); checkResult(2386, 3328);
        nextCycle(410); checkResult(2391, 3324);
        nextCycle(411); checkResult(2396, 3321);
        nextCycle(412); checkResult(2401, 3317);
        nextCycle(413); checkResult(2406, 3313);
        nextCycle(414); checkResult(2412, 3310);
        nextCycle(415); checkResult(2417, 3306);
        nextCycle(416); checkResult(2422, 3302);
        nextCycle(417); checkResult(2427, 3298);
        nextCycle(418); checkResult(2432, 3295);
        nextCycle(419); checkResult(2437, 3291);
        nextCycle(420); checkResult(2442, 3287);
        nextCycle(421); checkResult(2447, 3284);
        nextCycle(422); checkResult(2452, 3280);
        nextCycle(423); checkResult(2457, 3276);
        nextCycle(424); checkResult(2462, 3272);
        nextCycle(425); checkResult(2467, 3268);
        nextCycle(426); checkResult(2472, 3265);
        nextCycle(427); checkResult(2477, 3261);
        nextCycle(428); checkResult(2482, 3257);
        nextCycle(429); checkResult(2487, 3253);
        nextCycle(430); checkResult(2492, 3249);
        nextCycle(431); checkResult(2497, 3246);
        nextCycle(432); checkResult(2502, 3242);
        nextCycle(433); checkResult(2507, 3238);
        nextCycle(434); checkResult(2512, 3234);
        nextCycle(435); checkResult(2517, 3230);
        nextCycle(436); checkResult(2522, 3226);
        nextCycle(437); checkResult(2527, 3222);
        nextCycle(438); checkResult(2532, 3219);
        nextCycle(439); checkResult(2537, 3215);
        nextCycle(440); checkResult(2542, 3211);
        nextCycle(441); checkResult(2547, 3207);
        nextCycle(442); checkResult(2551, 3203);
        nextCycle(443); checkResult(2556, 3199);
        nextCycle(444); checkResult(2561, 3195);
        nextCycle(445); checkResult(2566, 3191);
        nextCycle(446); checkResult(2571, 3187);
        nextCycle(447); checkResult(2576, 3183);
        nextCycle(448); checkResult(2581, 3179);
        nextCycle(449); checkResult(2586, 3175);
        nextCycle(450); checkResult(2591, 3171);
        nextCycle(451); checkResult(2595, 3167);
        nextCycle(452); checkResult(2600, 3163);
        nextCycle(453); checkResult(2605, 3159);
        nextCycle(454); checkResult(2610, 3155);
        nextCycle(455); checkResult(2615, 3151);
        nextCycle(456); checkResult(2620, 3147);
        nextCycle(457); checkResult(2624, 3143);
        nextCycle(458); checkResult(2629, 3139);
        nextCycle(459); checkResult(2634, 3135);
        nextCycle(460); checkResult(2639, 3131);
        nextCycle(461); checkResult(2644, 3127);
        nextCycle(462); checkResult(2648, 3123);
        nextCycle(463); checkResult(2653, 3119);
        nextCycle(464); checkResult(2658, 3115);
        nextCycle(465); checkResult(2663, 3111);
        nextCycle(466); checkResult(2668, 3107);
        nextCycle(467); checkResult(2672, 3103);
        nextCycle(468); checkResult(2677, 3099);
        nextCycle(469); checkResult(2682, 3095);
        nextCycle(470); checkResult(2687, 3090);
        nextCycle(471); checkResult(2691, 3086);
        nextCycle(472); checkResult(2696, 3082);
        nextCycle(473); checkResult(2701, 3078);
        nextCycle(474); checkResult(2706, 3074);
        nextCycle(475); checkResult(2710, 3070);
        nextCycle(476); checkResult(2715, 3066);
        nextCycle(477); checkResult(2720, 3061);
        nextCycle(478); checkResult(2724, 3057);
        nextCycle(479); checkResult(2729, 3053);
        nextCycle(480); checkResult(2734, 3049);
        nextCycle(481); checkResult(2738, 3045);
        nextCycle(482); checkResult(2743, 3041);
        nextCycle(483); checkResult(2748, 3036);
        nextCycle(484); checkResult(2752, 3032);
        nextCycle(485); checkResult(2757, 3028);
        nextCycle(486); checkResult(2762, 3024);
        nextCycle(487); checkResult(2766, 3019);
        nextCycle(488); checkResult(2771, 3015);
        nextCycle(489); checkResult(2776, 3011);
        nextCycle(490); checkResult(2780, 3007);
        nextCycle(491); checkResult(2785, 3002);
        nextCycle(492); checkResult(2789, 2998);
        nextCycle(493); checkResult(2794, 2994);
        nextCycle(494); checkResult(2799, 2990);
        nextCycle(495); checkResult(2803, 2985);
        nextCycle(496); checkResult(2808, 2981);
        nextCycle(497); checkResult(2812, 2977);
        nextCycle(498); checkResult(2817, 2972);
        nextCycle(499); checkResult(2821, 2968);
        nextCycle(500); checkResult(2826, 2964);
        nextCycle(501); checkResult(2830, 2959);
        nextCycle(502); checkResult(2835, 2955);
        nextCycle(503); checkResult(2840, 2951);
        nextCycle(504); checkResult(2844, 2946);
        nextCycle(505); checkResult(2849, 2942);
        nextCycle(506); checkResult(2853, 2937);
        nextCycle(507); checkResult(2858, 2933);
        nextCycle(508); checkResult(2862, 2929);
        nextCycle(509); checkResult(2867, 2924);
        nextCycle(510); checkResult(2871, 2920);
        nextCycle(511); checkResult(2876, 2916);
        nextCycle(512); checkResult(2880, 2911);
        nextCycle(513); checkResult(2884, 2907);
        nextCycle(514); checkResult(2889, 2902);
        nextCycle(515); checkResult(2893, 2898);
        nextCycle(516); checkResult(2898, 2893);
        nextCycle(517); checkResult(2902, 2889);
        nextCycle(518); checkResult(2907, 2884);
        nextCycle(519); checkResult(2911, 2880);
        nextCycle(520); checkResult(2916, 2876);
        nextCycle(521); checkResult(2920, 2871);
        nextCycle(522); checkResult(2924, 2867);
        nextCycle(523); checkResult(2929, 2862);
        nextCycle(524); checkResult(2933, 2858);
        nextCycle(525); checkResult(2937, 2853);
        nextCycle(526); checkResult(2942, 2849);
        nextCycle(527); checkResult(2946, 2844);
        nextCycle(528); checkResult(2951, 2840);
        nextCycle(529); checkResult(2955, 2835);
        nextCycle(530); checkResult(2959, 2830);
        nextCycle(531); checkResult(2964, 2826);
        nextCycle(532); checkResult(2968, 2821);
        nextCycle(533); checkResult(2972, 2817);
        nextCycle(534); checkResult(2977, 2812);
        nextCycle(535); checkResult(2981, 2808);
        nextCycle(536); checkResult(2985, 2803);
        nextCycle(537); checkResult(2990, 2799);
        nextCycle(538); checkResult(2994, 2794);
        nextCycle(539); checkResult(2998, 2789);
        nextCycle(540); checkResult(3002, 2785);
        nextCycle(541); checkResult(3007, 2780);
        nextCycle(542); checkResult(3011, 2776);
        nextCycle(543); checkResult(3015, 2771);
        nextCycle(544); checkResult(3019, 2766);
        nextCycle(545); checkResult(3024, 2762);
        nextCycle(546); checkResult(3028, 2757);
        nextCycle(547); checkResult(3032, 2752);
        nextCycle(548); checkResult(3036, 2748);
        nextCycle(549); checkResult(3041, 2743);
        nextCycle(550); checkResult(3045, 2738);
        nextCycle(551); checkResult(3049, 2734);
        nextCycle(552); checkResult(3053, 2729);
        nextCycle(553); checkResult(3057, 2724);
        nextCycle(554); checkResult(3061, 2720);
        nextCycle(555); checkResult(3066, 2715);
        nextCycle(556); checkResult(3070, 2710);
        nextCycle(557); checkResult(3074, 2706);
        nextCycle(558); checkResult(3078, 2701);
        nextCycle(559); checkResult(3082, 2696);
        nextCycle(560); checkResult(3086, 2691);
        nextCycle(561); checkResult(3090, 2687);
        nextCycle(562); checkResult(3095, 2682);
        nextCycle(563); checkResult(3099, 2677);
        nextCycle(564); checkResult(3103, 2672);
        nextCycle(565); checkResult(3107, 2668);
        nextCycle(566); checkResult(3111, 2663);
        nextCycle(567); checkResult(3115, 2658);
        nextCycle(568); checkResult(3119, 2653);
        nextCycle(569); checkResult(3123, 2648);
        nextCycle(570); checkResult(3127, 2644);
        nextCycle(571); checkResult(3131, 2639);
        nextCycle(572); checkResult(3135, 2634);
        nextCycle(573); checkResult(3139, 2629);
        nextCycle(574); checkResult(3143, 2624);
        nextCycle(575); checkResult(3147, 2620);
        nextCycle(576); checkResult(3151, 2615);
        nextCycle(577); checkResult(3155, 2610);
        nextCycle(578); checkResult(3159, 2605);
        nextCycle(579); checkResult(3163, 2600);
        nextCycle(580); checkResult(3167, 2595);
        nextCycle(581); checkResult(3171, 2591);
        nextCycle(582); checkResult(3175, 2586);
        nextCycle(583); checkResult(3179, 2581);
        nextCycle(584); checkResult(3183, 2576);
        nextCycle(585); checkResult(3187, 2571);
        nextCycle(586); checkResult(3191, 2566);
        nextCycle(587); checkResult(3195, 2561);
        nextCycle(588); checkResult(3199, 2556);
        nextCycle(589); checkResult(3203, 2551);
        nextCycle(590); checkResult(3207, 2547);
        nextCycle(591); checkResult(3211, 2542);
        nextCycle(592); checkResult(3215, 2537);
        nextCycle(593); checkResult(3219, 2532);
        nextCycle(594); checkResult(3222, 2527);
        nextCycle(595); checkResult(3226, 2522);
        nextCycle(596); checkResult(3230, 2517);
        nextCycle(597); checkResult(3234, 2512);
        nextCycle(598); checkResult(3238, 2507);
        nextCycle(599); checkResult(3242, 2502);
        nextCycle(600); checkResult(3246, 2497);
        nextCycle(601); checkResult(3249, 2492);
        nextCycle(602); checkResult(3253, 2487);
        nextCycle(603); checkResult(3257, 2482);
        nextCycle(604); checkResult(3261, 2477);
        nextCycle(605); checkResult(3265, 2472);
        nextCycle(606); checkResult(3268, 2467);
        nextCycle(607); checkResult(3272, 2462);
        nextCycle(608); checkResult(3276, 2457);
        nextCycle(609); checkResult(3280, 2452);
        nextCycle(610); checkResult(3284, 2447);
        nextCycle(611); checkResult(3287, 2442);
        nextCycle(612); checkResult(3291, 2437);
        nextCycle(613); checkResult(3295, 2432);
        nextCycle(614); checkResult(3298, 2427);
        nextCycle(615); checkResult(3302, 2422);
        nextCycle(616); checkResult(3306, 2417);
        nextCycle(617); checkResult(3310, 2412);
        nextCycle(618); checkResult(3313, 2406);
        nextCycle(619); checkResult(3317, 2401);
        nextCycle(620); checkResult(3321, 2396);
        nextCycle(621); checkResult(3324, 2391);
        nextCycle(622); checkResult(3328, 2386);
        nextCycle(623); checkResult(3332, 2381);
        nextCycle(624); checkResult(3335, 2376);
        nextCycle(625); checkResult(3339, 2371);
        nextCycle(626); checkResult(3343, 2366);
        nextCycle(627); checkResult(3346, 2361);
        nextCycle(628); checkResult(3350, 2355);
        nextCycle(629); checkResult(3353, 2350);
        nextCycle(630); checkResult(3357, 2345);
        nextCycle(631); checkResult(3361, 2340);
        nextCycle(632); checkResult(3364, 2335);
        nextCycle(633); checkResult(3368, 2330);
        nextCycle(634); checkResult(3371, 2324);
        nextCycle(635); checkResult(3375, 2319);
        nextCycle(636); checkResult(3378, 2314);
        nextCycle(637); checkResult(3382, 2309);
        nextCycle(638); checkResult(3386, 2304);
        nextCycle(639); checkResult(3389, 2299);
        nextCycle(640); checkResult(3393, 2293);
        nextCycle(641); checkResult(3396, 2288);
        nextCycle(642); checkResult(3400, 2283);
        nextCycle(643); checkResult(3403, 2278);
        nextCycle(644); checkResult(3407, 2272);
        nextCycle(645); checkResult(3410, 2267);
        nextCycle(646); checkResult(3414, 2262);
        nextCycle(647); checkResult(3417, 2257);
        nextCycle(648); checkResult(3420, 2252);
        nextCycle(649); checkResult(3424, 2246);
        nextCycle(650); checkResult(3427, 2241);
        nextCycle(651); checkResult(3431, 2236);
        nextCycle(652); checkResult(3434, 2230);
        nextCycle(653); checkResult(3438, 2225);
        nextCycle(654); checkResult(3441, 2220);
        nextCycle(655); checkResult(3444, 2215);
        nextCycle(656); checkResult(3448, 2209);
        nextCycle(657); checkResult(3451, 2204);
        nextCycle(658); checkResult(3455, 2199);
        nextCycle(659); checkResult(3458, 2193);
        nextCycle(660); checkResult(3461, 2188);
        nextCycle(661); checkResult(3465, 2183);
        nextCycle(662); checkResult(3468, 2178);
        nextCycle(663); checkResult(3471, 2172);
        nextCycle(664); checkResult(3475, 2167);
        nextCycle(665); checkResult(3478, 2162);
        nextCycle(666); checkResult(3481, 2156);
        nextCycle(667); checkResult(3485, 2151);
        nextCycle(668); checkResult(3488, 2146);
        nextCycle(669); checkResult(3491, 2140);
        nextCycle(670); checkResult(3495, 2135);
        nextCycle(671); checkResult(3498, 2129);
        nextCycle(672); checkResult(3501, 2124);
        nextCycle(673); checkResult(3504, 2119);
        nextCycle(674); checkResult(3508, 2113);
        nextCycle(675); checkResult(3511, 2108);
        nextCycle(676); checkResult(3514, 2103);
        nextCycle(677); checkResult(3517, 2097);
        nextCycle(678); checkResult(3520, 2092);
        nextCycle(679); checkResult(3524, 2086);
        nextCycle(680); checkResult(3527, 2081);
        nextCycle(681); checkResult(3530, 2076);
        nextCycle(682); checkResult(3533, 2070);
        nextCycle(683); checkResult(3536, 2065);
        nextCycle(684); checkResult(3540, 2059);
        nextCycle(685); checkResult(3543, 2054);
        nextCycle(686); checkResult(3546, 2048);
        nextCycle(687); checkResult(3549, 2043);
        nextCycle(688); checkResult(3552, 2038);
        nextCycle(689); checkResult(3555, 2032);
        nextCycle(690); checkResult(3558, 2027);
        nextCycle(691); checkResult(3561, 2021);
        nextCycle(692); checkResult(3565, 2016);
        nextCycle(693); checkResult(3568, 2010);
        nextCycle(694); checkResult(3571, 2005);
        nextCycle(695); checkResult(3574, 1999);
        nextCycle(696); checkResult(3577, 1994);
        nextCycle(697); checkResult(3580, 1988);
        nextCycle(698); checkResult(3583, 1983);
        nextCycle(699); checkResult(3586, 1977);
        nextCycle(700); checkResult(3589, 1972);
        nextCycle(701); checkResult(3592, 1966);
        nextCycle(702); checkResult(3595, 1961);
        nextCycle(703); checkResult(3598, 1955);
        nextCycle(704); checkResult(3601, 1950);
        nextCycle(705); checkResult(3604, 1944);
        nextCycle(706); checkResult(3607, 1939);
        nextCycle(707); checkResult(3610, 1933);
        nextCycle(708); checkResult(3613, 1928);
        nextCycle(709); checkResult(3616, 1922);
        nextCycle(710); checkResult(3619, 1917);
        nextCycle(711); checkResult(3622, 1911);
        nextCycle(712); checkResult(3625, 1905);
        nextCycle(713); checkResult(3628, 1900);
        nextCycle(714); checkResult(3631, 1894);
        nextCycle(715); checkResult(3633, 1889);
        nextCycle(716); checkResult(3636, 1883);
        nextCycle(717); checkResult(3639, 1878);
        nextCycle(718); checkResult(3642, 1872);
        nextCycle(719); checkResult(3645, 1866);
        nextCycle(720); checkResult(3648, 1861);
        nextCycle(721); checkResult(3651, 1855);
        nextCycle(722); checkResult(3654, 1850);
        nextCycle(723); checkResult(3656, 1844);
        nextCycle(724); checkResult(3659, 1838);
        nextCycle(725); checkResult(3662, 1833);
        nextCycle(726); checkResult(3665, 1827);
        nextCycle(727); checkResult(3668, 1821);
        nextCycle(728); checkResult(3670, 1816);
        nextCycle(729); checkResult(3673, 1810);
        nextCycle(730); checkResult(3676, 1805);
        nextCycle(731); checkResult(3679, 1799);
        nextCycle(732); checkResult(3681, 1793);
        nextCycle(733); checkResult(3684, 1788);
        nextCycle(734); checkResult(3687, 1782);
        nextCycle(735); checkResult(3690, 1776);
        nextCycle(736); checkResult(3692, 1771);
        nextCycle(737); checkResult(3695, 1765);
        nextCycle(738); checkResult(3698, 1759);
        nextCycle(739); checkResult(3700, 1754);
        nextCycle(740); checkResult(3703, 1748);
        nextCycle(741); checkResult(3706, 1742);
        nextCycle(742); checkResult(3709, 1737);
        nextCycle(743); checkResult(3711, 1731);
        nextCycle(744); checkResult(3714, 1725);
        nextCycle(745); checkResult(3716, 1720);
        nextCycle(746); checkResult(3719, 1714);
        nextCycle(747); checkResult(3722, 1708);
        nextCycle(748); checkResult(3724, 1702);
        nextCycle(749); checkResult(3727, 1697);
        nextCycle(750); checkResult(3730, 1691);
        nextCycle(751); checkResult(3732, 1685);
        nextCycle(752); checkResult(3735, 1680);
        nextCycle(753); checkResult(3737, 1674);
        nextCycle(754); checkResult(3740, 1668);
        nextCycle(755); checkResult(3742, 1662);
        nextCycle(756); checkResult(3745, 1657);
        nextCycle(757); checkResult(3747, 1651);
        nextCycle(758); checkResult(3750, 1645);
        nextCycle(759); checkResult(3753, 1639);
        nextCycle(760); checkResult(3755, 1634);
        nextCycle(761); checkResult(3758, 1628);
        nextCycle(762); checkResult(3760, 1622);
        nextCycle(763); checkResult(3763, 1616);
        nextCycle(764); checkResult(3765, 1611);
        nextCycle(765); checkResult(3767, 1605);
        nextCycle(766); checkResult(3770, 1599);
        nextCycle(767); checkResult(3772, 1593);
        nextCycle(768); checkResult(3775, 1587);
        nextCycle(769); checkResult(3777, 1582);
        nextCycle(770); checkResult(3780, 1576);
        nextCycle(771); checkResult(3782, 1570);
        nextCycle(772); checkResult(3784, 1564);
        nextCycle(773); checkResult(3787, 1558);
        nextCycle(774); checkResult(3789, 1553);
        nextCycle(775); checkResult(3792, 1547);
        nextCycle(776); checkResult(3794, 1541);
        nextCycle(777); checkResult(3796, 1535);
        nextCycle(778); checkResult(3799, 1529);
        nextCycle(779); checkResult(3801, 1523);
        nextCycle(780); checkResult(3803, 1518);
        nextCycle(781); checkResult(3806, 1512);
        nextCycle(782); checkResult(3808, 1506);
        nextCycle(783); checkResult(3810, 1500);
        nextCycle(784); checkResult(3813, 1494);
        nextCycle(785); checkResult(3815, 1488);
        nextCycle(786); checkResult(3817, 1483);
        nextCycle(787); checkResult(3819, 1477);
        nextCycle(788); checkResult(3822, 1471);
        nextCycle(789); checkResult(3824, 1465);
        nextCycle(790); checkResult(3826, 1459);
        nextCycle(791); checkResult(3828, 1453);
        nextCycle(792); checkResult(3831, 1447);
        nextCycle(793); checkResult(3833, 1441);
        nextCycle(794); checkResult(3835, 1436);
        nextCycle(795); checkResult(3837, 1430);
        nextCycle(796); checkResult(3839, 1424);
        nextCycle(797); checkResult(3842, 1418);
        nextCycle(798); checkResult(3844, 1412);
        nextCycle(799); checkResult(3846, 1406);
        nextCycle(800); checkResult(3848, 1400);
        nextCycle(801); checkResult(3850, 1394);
        nextCycle(802); checkResult(3852, 1388);
        nextCycle(803); checkResult(3855, 1383);
        nextCycle(804); checkResult(3857, 1377);
        nextCycle(805); checkResult(3859, 1371);
        nextCycle(806); checkResult(3861, 1365);
        nextCycle(807); checkResult(3863, 1359);
        nextCycle(808); checkResult(3865, 1353);
        nextCycle(809); checkResult(3867, 1347);
        nextCycle(810); checkResult(3869, 1341);
        nextCycle(811); checkResult(3871, 1335);
        nextCycle(812); checkResult(3873, 1329);
        nextCycle(813); checkResult(3875, 1323);
        nextCycle(814); checkResult(3877, 1317);
        nextCycle(815); checkResult(3879, 1311);
        nextCycle(816); checkResult(3881, 1305);
        nextCycle(817); checkResult(3883, 1299);
        nextCycle(818); checkResult(3885, 1293);
        nextCycle(819); checkResult(3887, 1288);
        nextCycle(820); checkResult(3889, 1282);
        nextCycle(821); checkResult(3891, 1276);
        nextCycle(822); checkResult(3893, 1270);
        nextCycle(823); checkResult(3895, 1264);
        nextCycle(824); checkResult(3897, 1258);
        nextCycle(825); checkResult(3899, 1252);
        nextCycle(826); checkResult(3901, 1246);
        nextCycle(827); checkResult(3903, 1240);
        nextCycle(828); checkResult(3905, 1234);
        nextCycle(829); checkResult(3907, 1228);
        nextCycle(830); checkResult(3909, 1222);
        nextCycle(831); checkResult(3910, 1216);
        nextCycle(832); checkResult(3912, 1210);
        nextCycle(833); checkResult(3914, 1204);
        nextCycle(834); checkResult(3916, 1198);
        nextCycle(835); checkResult(3918, 1192);
        nextCycle(836); checkResult(3920, 1186);
        nextCycle(837); checkResult(3921, 1180);
        nextCycle(838); checkResult(3923, 1174);
        nextCycle(839); checkResult(3925, 1168);
        nextCycle(840); checkResult(3927, 1162);
        nextCycle(841); checkResult(3929, 1156);
        nextCycle(842); checkResult(3930, 1150);
        nextCycle(843); checkResult(3932, 1144);
        nextCycle(844); checkResult(3934, 1138);
        nextCycle(845); checkResult(3936, 1131);
        nextCycle(846); checkResult(3937, 1125);
        nextCycle(847); checkResult(3939, 1119);
        nextCycle(848); checkResult(3941, 1113);
        nextCycle(849); checkResult(3942, 1107);
        nextCycle(850); checkResult(3944, 1101);
        nextCycle(851); checkResult(3946, 1095);
        nextCycle(852); checkResult(3947, 1089);
        nextCycle(853); checkResult(3949, 1083);
        nextCycle(854); checkResult(3951, 1077);
        nextCycle(855); checkResult(3952, 1071);
        nextCycle(856); checkResult(3954, 1065);
        nextCycle(857); checkResult(3956, 1059);
        nextCycle(858); checkResult(3957, 1053);
        nextCycle(859); checkResult(3959, 1047);
        nextCycle(860); checkResult(3961, 1041);
        nextCycle(861); checkResult(3962, 1035);
        nextCycle(862); checkResult(3964, 1028);
        nextCycle(863); checkResult(3965, 1022);
        nextCycle(864); checkResult(3967, 1016);
        nextCycle(865); checkResult(3968, 1010);
        nextCycle(866); checkResult(3970, 1004);
        nextCycle(867); checkResult(3972, 998);
        nextCycle(868); checkResult(3973, 992);
        nextCycle(869); checkResult(3975, 986);
        nextCycle(870); checkResult(3976, 980);
        nextCycle(871); checkResult(3978, 974);
        nextCycle(872); checkResult(3979, 968);
        nextCycle(873); checkResult(3981, 961);
        nextCycle(874); checkResult(3982, 955);
        nextCycle(875); checkResult(3983, 949);
        nextCycle(876); checkResult(3985, 943);
        nextCycle(877); checkResult(3986, 937);
        nextCycle(878); checkResult(3988, 931);
        nextCycle(879); checkResult(3989, 925);
        nextCycle(880); checkResult(3991, 919);
        nextCycle(881); checkResult(3992, 913);
        nextCycle(882); checkResult(3993, 906);
        nextCycle(883); checkResult(3995, 900);
        nextCycle(884); checkResult(3996, 894);
        nextCycle(885); checkResult(3998, 888);
        nextCycle(886); checkResult(3999, 882);
        nextCycle(887); checkResult(4000, 876);
        nextCycle(888); checkResult(4002, 870);
        nextCycle(889); checkResult(4003, 863);
        nextCycle(890); checkResult(4004, 857);
        nextCycle(891); checkResult(4006, 851);
        nextCycle(892); checkResult(4007, 845);
        nextCycle(893); checkResult(4008, 839);
        nextCycle(894); checkResult(4009, 833);
        nextCycle(895); checkResult(4011, 827);
        nextCycle(896); checkResult(4012, 820);
        nextCycle(897); checkResult(4013, 814);
        nextCycle(898); checkResult(4014, 808);
        nextCycle(899); checkResult(4016, 802);
        nextCycle(900); checkResult(4017, 796);
        nextCycle(901); checkResult(4018, 790);
        nextCycle(902); checkResult(4019, 783);
        nextCycle(903); checkResult(4021, 777);
        nextCycle(904); checkResult(4022, 771);
        nextCycle(905); checkResult(4023, 765);
        nextCycle(906); checkResult(4024, 759);
        nextCycle(907); checkResult(4025, 753);
        nextCycle(908); checkResult(4026, 746);
        nextCycle(909); checkResult(4028, 740);
        nextCycle(910); checkResult(4029, 734);
        nextCycle(911); checkResult(4030, 728);
        nextCycle(912); checkResult(4031, 722);
        nextCycle(913); checkResult(4032, 716);
        nextCycle(914); checkResult(4033, 709);
        nextCycle(915); checkResult(4034, 703);
        nextCycle(916); checkResult(4035, 697);
        nextCycle(917); checkResult(4036, 691);
        nextCycle(918); checkResult(4037, 685);
        nextCycle(919); checkResult(4038, 678);
        nextCycle(920); checkResult(4039, 672);
        nextCycle(921); checkResult(4040, 666);
        nextCycle(922); checkResult(4041, 660);
        nextCycle(923); checkResult(4042, 654);
        nextCycle(924); checkResult(4043, 647);
        nextCycle(925); checkResult(4044, 641);
        nextCycle(926); checkResult(4045, 635);
        nextCycle(927); checkResult(4046, 629);
        nextCycle(928); checkResult(4047, 623);
        nextCycle(929); checkResult(4048, 616);
        nextCycle(930); checkResult(4049, 610);
        nextCycle(931); checkResult(4050, 604);
        nextCycle(932); checkResult(4051, 598);
        nextCycle(933); checkResult(4052, 592);
        nextCycle(934); checkResult(4053, 585);
        nextCycle(935); checkResult(4054, 579);
        nextCycle(936); checkResult(4055, 573);
        nextCycle(937); checkResult(4056, 567);
        nextCycle(938); checkResult(4056, 560);
        nextCycle(939); checkResult(4057, 554);
        nextCycle(940); checkResult(4058, 548);
        nextCycle(941); checkResult(4059, 542);
        nextCycle(942); checkResult(4060, 536);
        nextCycle(943); checkResult(4061, 529);
        nextCycle(944); checkResult(4061, 523);
        nextCycle(945); checkResult(4062, 517);
        nextCycle(946); checkResult(4063, 511);
        nextCycle(947); checkResult(4064, 504);
        nextCycle(948); checkResult(4065, 498);
        nextCycle(949); checkResult(4065, 492);
        nextCycle(950); checkResult(4066, 486);
        nextCycle(951); checkResult(4067, 479);
        nextCycle(952); checkResult(4068, 473);
        nextCycle(953); checkResult(4068, 467);
        nextCycle(954); checkResult(4069, 461);
        nextCycle(955); checkResult(4070, 454);
        nextCycle(956); checkResult(4070, 448);
        nextCycle(957); checkResult(4071, 442);
        nextCycle(958); checkResult(4072, 436);
        nextCycle(959); checkResult(4072, 430);
        nextCycle(960); checkResult(4073, 423);
        nextCycle(961); checkResult(4074, 417);
        nextCycle(962); checkResult(4074, 411);
        nextCycle(963); checkResult(4075, 405);
        nextCycle(964); checkResult(4076, 398);
        nextCycle(965); checkResult(4076, 392);
        nextCycle(966); checkResult(4077, 386);
        nextCycle(967); checkResult(4077, 379);
        nextCycle(968); checkResult(4078, 373);
        nextCycle(969); checkResult(4079, 367);
        nextCycle(970); checkResult(4079, 361);
        nextCycle(971); checkResult(4080, 354);
        nextCycle(972); checkResult(4080, 348);
        nextCycle(973); checkResult(4081, 342);
        nextCycle(974); checkResult(4081, 336);
        nextCycle(975); checkResult(4082, 329);
        nextCycle(976); checkResult(4082, 323);
        nextCycle(977); checkResult(4083, 317);
        nextCycle(978); checkResult(4083, 311);
        nextCycle(979); checkResult(4084, 304);
        nextCycle(980); checkResult(4084, 298);
        nextCycle(981); checkResult(4085, 292);
        nextCycle(982); checkResult(4085, 286);
        nextCycle(983); checkResult(4085, 279);
        nextCycle(984); checkResult(4086, 273);
        nextCycle(985); checkResult(4086, 267);
        nextCycle(986); checkResult(4087, 261);
        nextCycle(987); checkResult(4087, 254);
        nextCycle(988); checkResult(4087, 248);
        nextCycle(989); checkResult(4088, 242);
        nextCycle(990); checkResult(4088, 235);
        nextCycle(991); checkResult(4089, 229);
        nextCycle(992); checkResult(4089, 223);
        nextCycle(993); checkResult(4089, 217);
        nextCycle(994); checkResult(4090, 210);
        nextCycle(995); checkResult(4090, 204);
        nextCycle(996); checkResult(4090, 198);
        nextCycle(997); checkResult(4091, 192);
        nextCycle(998); checkResult(4091, 185);
        nextCycle(999); checkResult(4091, 179);
        nextCycle(1000); checkResult(4091, 173);
        nextCycle(1001); checkResult(4092, 166);
        nextCycle(1002); checkResult(4092, 160);
        nextCycle(1003); checkResult(4092, 154);
        nextCycle(1004); checkResult(4092, 148);
        nextCycle(1005); checkResult(4093, 141);
        nextCycle(1006); checkResult(4093, 135);
        nextCycle(1007); checkResult(4093, 129);
        nextCycle(1008); checkResult(4093, 122);
        nextCycle(1009); checkResult(4093, 116);
        nextCycle(1010); checkResult(4094, 110);
        nextCycle(1011); checkResult(4094, 104);
        nextCycle(1012); checkResult(4094, 97);
        nextCycle(1013); checkResult(4094, 91);
        nextCycle(1014); checkResult(4094, 85);
        nextCycle(1015); checkResult(4094, 79);
        nextCycle(1016); checkResult(4094, 72);
        nextCycle(1017); checkResult(4094, 66);
        nextCycle(1018); checkResult(4095, 60);
        nextCycle(1019); checkResult(4095, 53);
        nextCycle(1020); checkResult(4095, 47);
        nextCycle(1021); checkResult(4095, 41);
        nextCycle(1022); checkResult(4095, 35);
        nextCycle(1023); checkResult(4095, 28);
        nextCycle(1024); checkResult(4095, 22);
        nextCycle(1025); checkResult(4095, 16);
        nextCycle(1026); checkResult(4095, 9);
        nextCycle(1027); checkResult(4095, 3);
        nextCycle(1028); checkResult(4095, -3);
        nextCycle(1029); checkResult(4095, -9);
        nextCycle(1030); checkResult(4095, -16);
        nextCycle(1031); checkResult(4095, -22);
        nextCycle(1032); checkResult(4095, -28);
        nextCycle(1033); checkResult(4095, -35);
        nextCycle(1034); checkResult(4095, -41);
        nextCycle(1035); checkResult(4095, -47);
        nextCycle(1036); checkResult(4095, -53);
        nextCycle(1037); checkResult(4095, -60);
        nextCycle(1038); checkResult(4094, -66);
        nextCycle(1039); checkResult(4094, -72);
        nextCycle(1040); checkResult(4094, -79);
        nextCycle(1041); checkResult(4094, -85);
        nextCycle(1042); checkResult(4094, -91);
        nextCycle(1043); checkResult(4094, -97);
        nextCycle(1044); checkResult(4094, -104);
        nextCycle(1045); checkResult(4094, -110);
        nextCycle(1046); checkResult(4093, -116);
        nextCycle(1047); checkResult(4093, -122);
        nextCycle(1048); checkResult(4093, -129);
        nextCycle(1049); checkResult(4093, -135);
        nextCycle(1050); checkResult(4093, -141);
        nextCycle(1051); checkResult(4092, -148);
        nextCycle(1052); checkResult(4092, -154);
        nextCycle(1053); checkResult(4092, -160);
        nextCycle(1054); checkResult(4092, -166);
        nextCycle(1055); checkResult(4091, -173);
        nextCycle(1056); checkResult(4091, -179);
        nextCycle(1057); checkResult(4091, -185);
        nextCycle(1058); checkResult(4091, -192);
        nextCycle(1059); checkResult(4090, -198);
        nextCycle(1060); checkResult(4090, -204);
        nextCycle(1061); checkResult(4090, -210);
        nextCycle(1062); checkResult(4089, -217);
        nextCycle(1063); checkResult(4089, -223);
        nextCycle(1064); checkResult(4089, -229);
        nextCycle(1065); checkResult(4088, -235);
        nextCycle(1066); checkResult(4088, -242);
        nextCycle(1067); checkResult(4087, -248);
        nextCycle(1068); checkResult(4087, -254);
        nextCycle(1069); checkResult(4087, -261);
        nextCycle(1070); checkResult(4086, -267);
        nextCycle(1071); checkResult(4086, -273);
        nextCycle(1072); checkResult(4085, -279);
        nextCycle(1073); checkResult(4085, -286);
        nextCycle(1074); checkResult(4085, -292);
        nextCycle(1075); checkResult(4084, -298);
        nextCycle(1076); checkResult(4084, -304);
        nextCycle(1077); checkResult(4083, -311);
        nextCycle(1078); checkResult(4083, -317);
        nextCycle(1079); checkResult(4082, -323);
        nextCycle(1080); checkResult(4082, -329);
        nextCycle(1081); checkResult(4081, -336);
        nextCycle(1082); checkResult(4081, -342);
        nextCycle(1083); checkResult(4080, -348);
        nextCycle(1084); checkResult(4080, -354);
        nextCycle(1085); checkResult(4079, -361);
        nextCycle(1086); checkResult(4079, -367);
        nextCycle(1087); checkResult(4078, -373);
        nextCycle(1088); checkResult(4077, -379);
        nextCycle(1089); checkResult(4077, -386);
        nextCycle(1090); checkResult(4076, -392);
        nextCycle(1091); checkResult(4076, -398);
        nextCycle(1092); checkResult(4075, -405);
        nextCycle(1093); checkResult(4074, -411);
        nextCycle(1094); checkResult(4074, -417);
        nextCycle(1095); checkResult(4073, -423);
        nextCycle(1096); checkResult(4072, -430);
        nextCycle(1097); checkResult(4072, -436);
        nextCycle(1098); checkResult(4071, -442);
        nextCycle(1099); checkResult(4070, -448);
        nextCycle(1100); checkResult(4070, -454);
        nextCycle(1101); checkResult(4069, -461);
        nextCycle(1102); checkResult(4068, -467);
        nextCycle(1103); checkResult(4068, -473);
        nextCycle(1104); checkResult(4067, -479);
        nextCycle(1105); checkResult(4066, -486);
        nextCycle(1106); checkResult(4065, -492);
        nextCycle(1107); checkResult(4065, -498);
        nextCycle(1108); checkResult(4064, -504);
        nextCycle(1109); checkResult(4063, -511);
        nextCycle(1110); checkResult(4062, -517);
        nextCycle(1111); checkResult(4061, -523);
        nextCycle(1112); checkResult(4061, -529);
        nextCycle(1113); checkResult(4060, -536);
        nextCycle(1114); checkResult(4059, -542);
        nextCycle(1115); checkResult(4058, -548);
        nextCycle(1116); checkResult(4057, -554);
        nextCycle(1117); checkResult(4056, -560);
        nextCycle(1118); checkResult(4056, -567);
        nextCycle(1119); checkResult(4055, -573);
        nextCycle(1120); checkResult(4054, -579);
        nextCycle(1121); checkResult(4053, -585);
        nextCycle(1122); checkResult(4052, -592);
        nextCycle(1123); checkResult(4051, -598);
        nextCycle(1124); checkResult(4050, -604);
        nextCycle(1125); checkResult(4049, -610);
        nextCycle(1126); checkResult(4048, -616);
        nextCycle(1127); checkResult(4047, -623);
        nextCycle(1128); checkResult(4046, -629);
        nextCycle(1129); checkResult(4045, -635);
        nextCycle(1130); checkResult(4044, -641);
        nextCycle(1131); checkResult(4043, -647);
        nextCycle(1132); checkResult(4042, -654);
        nextCycle(1133); checkResult(4041, -660);
        nextCycle(1134); checkResult(4040, -666);
        nextCycle(1135); checkResult(4039, -672);
        nextCycle(1136); checkResult(4038, -678);
        nextCycle(1137); checkResult(4037, -685);
        nextCycle(1138); checkResult(4036, -691);
        nextCycle(1139); checkResult(4035, -697);
        nextCycle(1140); checkResult(4034, -703);
        nextCycle(1141); checkResult(4033, -709);
        nextCycle(1142); checkResult(4032, -716);
        nextCycle(1143); checkResult(4031, -722);
        nextCycle(1144); checkResult(4030, -728);
        nextCycle(1145); checkResult(4029, -734);
        nextCycle(1146); checkResult(4028, -740);
        nextCycle(1147); checkResult(4026, -746);
        nextCycle(1148); checkResult(4025, -753);
        nextCycle(1149); checkResult(4024, -759);
        nextCycle(1150); checkResult(4023, -765);
        nextCycle(1151); checkResult(4022, -771);
        nextCycle(1152); checkResult(4021, -777);
        nextCycle(1153); checkResult(4019, -783);
        nextCycle(1154); checkResult(4018, -790);
        nextCycle(1155); checkResult(4017, -796);
        nextCycle(1156); checkResult(4016, -802);
        nextCycle(1157); checkResult(4014, -808);
        nextCycle(1158); checkResult(4013, -814);
        nextCycle(1159); checkResult(4012, -820);
        nextCycle(1160); checkResult(4011, -827);
        nextCycle(1161); checkResult(4009, -833);
        nextCycle(1162); checkResult(4008, -839);
        nextCycle(1163); checkResult(4007, -845);
        nextCycle(1164); checkResult(4006, -851);
        nextCycle(1165); checkResult(4004, -857);
        nextCycle(1166); checkResult(4003, -863);
        nextCycle(1167); checkResult(4002, -870);
        nextCycle(1168); checkResult(4000, -876);
        nextCycle(1169); checkResult(3999, -882);
        nextCycle(1170); checkResult(3998, -888);
        nextCycle(1171); checkResult(3996, -894);
        nextCycle(1172); checkResult(3995, -900);
        nextCycle(1173); checkResult(3993, -906);
        nextCycle(1174); checkResult(3992, -913);
        nextCycle(1175); checkResult(3991, -919);
        nextCycle(1176); checkResult(3989, -925);
        nextCycle(1177); checkResult(3988, -931);
        nextCycle(1178); checkResult(3986, -937);
        nextCycle(1179); checkResult(3985, -943);
        nextCycle(1180); checkResult(3983, -949);
        nextCycle(1181); checkResult(3982, -955);
        nextCycle(1182); checkResult(3981, -961);
        nextCycle(1183); checkResult(3979, -968);
        nextCycle(1184); checkResult(3978, -974);
        nextCycle(1185); checkResult(3976, -980);
        nextCycle(1186); checkResult(3975, -986);
        nextCycle(1187); checkResult(3973, -992);
        nextCycle(1188); checkResult(3972, -998);
        nextCycle(1189); checkResult(3970, -1004);
        nextCycle(1190); checkResult(3968, -1010);
        nextCycle(1191); checkResult(3967, -1016);
        nextCycle(1192); checkResult(3965, -1022);
        nextCycle(1193); checkResult(3964, -1028);
        nextCycle(1194); checkResult(3962, -1035);
        nextCycle(1195); checkResult(3961, -1041);
        nextCycle(1196); checkResult(3959, -1047);
        nextCycle(1197); checkResult(3957, -1053);
        nextCycle(1198); checkResult(3956, -1059);
        nextCycle(1199); checkResult(3954, -1065);
        nextCycle(1200); checkResult(3952, -1071);
        nextCycle(1201); checkResult(3951, -1077);
        nextCycle(1202); checkResult(3949, -1083);
        nextCycle(1203); checkResult(3947, -1089);
        nextCycle(1204); checkResult(3946, -1095);
        nextCycle(1205); checkResult(3944, -1101);
        nextCycle(1206); checkResult(3942, -1107);
        nextCycle(1207); checkResult(3941, -1113);
        nextCycle(1208); checkResult(3939, -1119);
        nextCycle(1209); checkResult(3937, -1125);
        nextCycle(1210); checkResult(3936, -1131);
        nextCycle(1211); checkResult(3934, -1138);
        nextCycle(1212); checkResult(3932, -1144);
        nextCycle(1213); checkResult(3930, -1150);
        nextCycle(1214); checkResult(3929, -1156);
        nextCycle(1215); checkResult(3927, -1162);
        nextCycle(1216); checkResult(3925, -1168);
        nextCycle(1217); checkResult(3923, -1174);
        nextCycle(1218); checkResult(3921, -1180);
        nextCycle(1219); checkResult(3920, -1186);
        nextCycle(1220); checkResult(3918, -1192);
        nextCycle(1221); checkResult(3916, -1198);
        nextCycle(1222); checkResult(3914, -1204);
        nextCycle(1223); checkResult(3912, -1210);
        nextCycle(1224); checkResult(3910, -1216);
        nextCycle(1225); checkResult(3909, -1222);
        nextCycle(1226); checkResult(3907, -1228);
        nextCycle(1227); checkResult(3905, -1234);
        nextCycle(1228); checkResult(3903, -1240);
        nextCycle(1229); checkResult(3901, -1246);
        nextCycle(1230); checkResult(3899, -1252);
        nextCycle(1231); checkResult(3897, -1258);
        nextCycle(1232); checkResult(3895, -1264);
        nextCycle(1233); checkResult(3893, -1270);
        nextCycle(1234); checkResult(3891, -1276);
        nextCycle(1235); checkResult(3889, -1282);
        nextCycle(1236); checkResult(3887, -1288);
        nextCycle(1237); checkResult(3885, -1293);
        nextCycle(1238); checkResult(3883, -1299);
        nextCycle(1239); checkResult(3881, -1305);
        nextCycle(1240); checkResult(3879, -1311);
        nextCycle(1241); checkResult(3877, -1317);
        nextCycle(1242); checkResult(3875, -1323);
        nextCycle(1243); checkResult(3873, -1329);
        nextCycle(1244); checkResult(3871, -1335);
        nextCycle(1245); checkResult(3869, -1341);
        nextCycle(1246); checkResult(3867, -1347);
        nextCycle(1247); checkResult(3865, -1353);
        nextCycle(1248); checkResult(3863, -1359);
        nextCycle(1249); checkResult(3861, -1365);
        nextCycle(1250); checkResult(3859, -1371);
        nextCycle(1251); checkResult(3857, -1377);
        nextCycle(1252); checkResult(3855, -1383);
        nextCycle(1253); checkResult(3852, -1388);
        nextCycle(1254); checkResult(3850, -1394);
        nextCycle(1255); checkResult(3848, -1400);
        nextCycle(1256); checkResult(3846, -1406);
        nextCycle(1257); checkResult(3844, -1412);
        nextCycle(1258); checkResult(3842, -1418);
        nextCycle(1259); checkResult(3839, -1424);
        nextCycle(1260); checkResult(3837, -1430);
        nextCycle(1261); checkResult(3835, -1436);
        nextCycle(1262); checkResult(3833, -1441);
        nextCycle(1263); checkResult(3831, -1447);
        nextCycle(1264); checkResult(3828, -1453);
        nextCycle(1265); checkResult(3826, -1459);
        nextCycle(1266); checkResult(3824, -1465);
        nextCycle(1267); checkResult(3822, -1471);
        nextCycle(1268); checkResult(3819, -1477);
        nextCycle(1269); checkResult(3817, -1483);
        nextCycle(1270); checkResult(3815, -1488);
        nextCycle(1271); checkResult(3813, -1494);
        nextCycle(1272); checkResult(3810, -1500);
        nextCycle(1273); checkResult(3808, -1506);
        nextCycle(1274); checkResult(3806, -1512);
        nextCycle(1275); checkResult(3803, -1518);
        nextCycle(1276); checkResult(3801, -1523);
        nextCycle(1277); checkResult(3799, -1529);
        nextCycle(1278); checkResult(3796, -1535);
        nextCycle(1279); checkResult(3794, -1541);
        nextCycle(1280); checkResult(3792, -1547);
        nextCycle(1281); checkResult(3789, -1553);
        nextCycle(1282); checkResult(3787, -1558);
        nextCycle(1283); checkResult(3784, -1564);
        nextCycle(1284); checkResult(3782, -1570);
        nextCycle(1285); checkResult(3780, -1576);
        nextCycle(1286); checkResult(3777, -1582);
        nextCycle(1287); checkResult(3775, -1587);
        nextCycle(1288); checkResult(3772, -1593);
        nextCycle(1289); checkResult(3770, -1599);
        nextCycle(1290); checkResult(3767, -1605);
        nextCycle(1291); checkResult(3765, -1611);
        nextCycle(1292); checkResult(3763, -1616);
        nextCycle(1293); checkResult(3760, -1622);
        nextCycle(1294); checkResult(3758, -1628);
        nextCycle(1295); checkResult(3755, -1634);
        nextCycle(1296); checkResult(3753, -1639);
        nextCycle(1297); checkResult(3750, -1645);
        nextCycle(1298); checkResult(3747, -1651);
        nextCycle(1299); checkResult(3745, -1657);
        nextCycle(1300); checkResult(3742, -1662);
        nextCycle(1301); checkResult(3740, -1668);
        nextCycle(1302); checkResult(3737, -1674);
        nextCycle(1303); checkResult(3735, -1680);
        nextCycle(1304); checkResult(3732, -1685);
        nextCycle(1305); checkResult(3730, -1691);
        nextCycle(1306); checkResult(3727, -1697);
        nextCycle(1307); checkResult(3724, -1702);
        nextCycle(1308); checkResult(3722, -1708);
        nextCycle(1309); checkResult(3719, -1714);
        nextCycle(1310); checkResult(3716, -1720);
        nextCycle(1311); checkResult(3714, -1725);
        nextCycle(1312); checkResult(3711, -1731);
        nextCycle(1313); checkResult(3709, -1737);
        nextCycle(1314); checkResult(3706, -1742);
        nextCycle(1315); checkResult(3703, -1748);
        nextCycle(1316); checkResult(3700, -1754);
        nextCycle(1317); checkResult(3698, -1759);
        nextCycle(1318); checkResult(3695, -1765);
        nextCycle(1319); checkResult(3692, -1771);
        nextCycle(1320); checkResult(3690, -1776);
        nextCycle(1321); checkResult(3687, -1782);
        nextCycle(1322); checkResult(3684, -1788);
        nextCycle(1323); checkResult(3681, -1793);
        nextCycle(1324); checkResult(3679, -1799);
        nextCycle(1325); checkResult(3676, -1805);
        nextCycle(1326); checkResult(3673, -1810);
        nextCycle(1327); checkResult(3670, -1816);
        nextCycle(1328); checkResult(3668, -1821);
        nextCycle(1329); checkResult(3665, -1827);
        nextCycle(1330); checkResult(3662, -1833);
        nextCycle(1331); checkResult(3659, -1838);
        nextCycle(1332); checkResult(3656, -1844);
        nextCycle(1333); checkResult(3654, -1850);
        nextCycle(1334); checkResult(3651, -1855);
        nextCycle(1335); checkResult(3648, -1861);
        nextCycle(1336); checkResult(3645, -1866);
        nextCycle(1337); checkResult(3642, -1872);
        nextCycle(1338); checkResult(3639, -1878);
        nextCycle(1339); checkResult(3636, -1883);
        nextCycle(1340); checkResult(3633, -1889);
        nextCycle(1341); checkResult(3631, -1894);
        nextCycle(1342); checkResult(3628, -1900);
        nextCycle(1343); checkResult(3625, -1905);
        nextCycle(1344); checkResult(3622, -1911);
        nextCycle(1345); checkResult(3619, -1917);
        nextCycle(1346); checkResult(3616, -1922);
        nextCycle(1347); checkResult(3613, -1928);
        nextCycle(1348); checkResult(3610, -1933);
        nextCycle(1349); checkResult(3607, -1939);
        nextCycle(1350); checkResult(3604, -1944);
        nextCycle(1351); checkResult(3601, -1950);
        nextCycle(1352); checkResult(3598, -1955);
        nextCycle(1353); checkResult(3595, -1961);
        nextCycle(1354); checkResult(3592, -1966);
        nextCycle(1355); checkResult(3589, -1972);
        nextCycle(1356); checkResult(3586, -1977);
        nextCycle(1357); checkResult(3583, -1983);
        nextCycle(1358); checkResult(3580, -1988);
        nextCycle(1359); checkResult(3577, -1994);
        nextCycle(1360); checkResult(3574, -1999);
        nextCycle(1361); checkResult(3571, -2005);
        nextCycle(1362); checkResult(3568, -2010);
        nextCycle(1363); checkResult(3565, -2016);
        nextCycle(1364); checkResult(3561, -2021);
        nextCycle(1365); checkResult(3558, -2027);
        nextCycle(1366); checkResult(3555, -2032);
        nextCycle(1367); checkResult(3552, -2038);
        nextCycle(1368); checkResult(3549, -2043);
        nextCycle(1369); checkResult(3546, -2048);
        nextCycle(1370); checkResult(3543, -2054);
        nextCycle(1371); checkResult(3540, -2059);
        nextCycle(1372); checkResult(3536, -2065);
        nextCycle(1373); checkResult(3533, -2070);
        nextCycle(1374); checkResult(3530, -2076);
        nextCycle(1375); checkResult(3527, -2081);
        nextCycle(1376); checkResult(3524, -2086);
        nextCycle(1377); checkResult(3520, -2092);
        nextCycle(1378); checkResult(3517, -2097);
        nextCycle(1379); checkResult(3514, -2103);
        nextCycle(1380); checkResult(3511, -2108);
        nextCycle(1381); checkResult(3508, -2113);
        nextCycle(1382); checkResult(3504, -2119);
        nextCycle(1383); checkResult(3501, -2124);
        nextCycle(1384); checkResult(3498, -2129);
        nextCycle(1385); checkResult(3495, -2135);
        nextCycle(1386); checkResult(3491, -2140);
        nextCycle(1387); checkResult(3488, -2146);
        nextCycle(1388); checkResult(3485, -2151);
        nextCycle(1389); checkResult(3481, -2156);
        nextCycle(1390); checkResult(3478, -2162);
        nextCycle(1391); checkResult(3475, -2167);
        nextCycle(1392); checkResult(3471, -2172);
        nextCycle(1393); checkResult(3468, -2178);
        nextCycle(1394); checkResult(3465, -2183);
        nextCycle(1395); checkResult(3461, -2188);
        nextCycle(1396); checkResult(3458, -2193);
        nextCycle(1397); checkResult(3455, -2199);
        nextCycle(1398); checkResult(3451, -2204);
        nextCycle(1399); checkResult(3448, -2209);
        nextCycle(1400); checkResult(3444, -2215);
        nextCycle(1401); checkResult(3441, -2220);
        nextCycle(1402); checkResult(3438, -2225);
        nextCycle(1403); checkResult(3434, -2230);
        nextCycle(1404); checkResult(3431, -2236);
        nextCycle(1405); checkResult(3427, -2241);
        nextCycle(1406); checkResult(3424, -2246);
        nextCycle(1407); checkResult(3420, -2252);
        nextCycle(1408); checkResult(3417, -2257);
        nextCycle(1409); checkResult(3414, -2262);
        nextCycle(1410); checkResult(3410, -2267);
        nextCycle(1411); checkResult(3407, -2272);
        nextCycle(1412); checkResult(3403, -2278);
        nextCycle(1413); checkResult(3400, -2283);
        nextCycle(1414); checkResult(3396, -2288);
        nextCycle(1415); checkResult(3393, -2293);
        nextCycle(1416); checkResult(3389, -2299);
        nextCycle(1417); checkResult(3386, -2304);
        nextCycle(1418); checkResult(3382, -2309);
        nextCycle(1419); checkResult(3378, -2314);
        nextCycle(1420); checkResult(3375, -2319);
        nextCycle(1421); checkResult(3371, -2324);
        nextCycle(1422); checkResult(3368, -2330);
        nextCycle(1423); checkResult(3364, -2335);
        nextCycle(1424); checkResult(3361, -2340);
        nextCycle(1425); checkResult(3357, -2345);
        nextCycle(1426); checkResult(3353, -2350);
        nextCycle(1427); checkResult(3350, -2355);
        nextCycle(1428); checkResult(3346, -2361);
        nextCycle(1429); checkResult(3343, -2366);
        nextCycle(1430); checkResult(3339, -2371);
        nextCycle(1431); checkResult(3335, -2376);
        nextCycle(1432); checkResult(3332, -2381);
        nextCycle(1433); checkResult(3328, -2386);
        nextCycle(1434); checkResult(3324, -2391);
        nextCycle(1435); checkResult(3321, -2396);
        nextCycle(1436); checkResult(3317, -2401);
        nextCycle(1437); checkResult(3313, -2406);
        nextCycle(1438); checkResult(3310, -2412);
        nextCycle(1439); checkResult(3306, -2417);
        nextCycle(1440); checkResult(3302, -2422);
        nextCycle(1441); checkResult(3298, -2427);
        nextCycle(1442); checkResult(3295, -2432);
        nextCycle(1443); checkResult(3291, -2437);
        nextCycle(1444); checkResult(3287, -2442);
        nextCycle(1445); checkResult(3284, -2447);
        nextCycle(1446); checkResult(3280, -2452);
        nextCycle(1447); checkResult(3276, -2457);
        nextCycle(1448); checkResult(3272, -2462);
        nextCycle(1449); checkResult(3268, -2467);
        nextCycle(1450); checkResult(3265, -2472);
        nextCycle(1451); checkResult(3261, -2477);
        nextCycle(1452); checkResult(3257, -2482);
        nextCycle(1453); checkResult(3253, -2487);
        nextCycle(1454); checkResult(3249, -2492);
        nextCycle(1455); checkResult(3246, -2497);
        nextCycle(1456); checkResult(3242, -2502);
        nextCycle(1457); checkResult(3238, -2507);
        nextCycle(1458); checkResult(3234, -2512);
        nextCycle(1459); checkResult(3230, -2517);
        nextCycle(1460); checkResult(3226, -2522);
        nextCycle(1461); checkResult(3222, -2527);
        nextCycle(1462); checkResult(3219, -2532);
        nextCycle(1463); checkResult(3215, -2537);
        nextCycle(1464); checkResult(3211, -2542);
        nextCycle(1465); checkResult(3207, -2547);
        nextCycle(1466); checkResult(3203, -2551);
        nextCycle(1467); checkResult(3199, -2556);
        nextCycle(1468); checkResult(3195, -2561);
        nextCycle(1469); checkResult(3191, -2566);
        nextCycle(1470); checkResult(3187, -2571);
        nextCycle(1471); checkResult(3183, -2576);
        nextCycle(1472); checkResult(3179, -2581);
        nextCycle(1473); checkResult(3175, -2586);
        nextCycle(1474); checkResult(3171, -2591);
        nextCycle(1475); checkResult(3167, -2595);
        nextCycle(1476); checkResult(3163, -2600);
        nextCycle(1477); checkResult(3159, -2605);
        nextCycle(1478); checkResult(3155, -2610);
        nextCycle(1479); checkResult(3151, -2615);
        nextCycle(1480); checkResult(3147, -2620);
        nextCycle(1481); checkResult(3143, -2624);
        nextCycle(1482); checkResult(3139, -2629);
        nextCycle(1483); checkResult(3135, -2634);
        nextCycle(1484); checkResult(3131, -2639);
        nextCycle(1485); checkResult(3127, -2644);
        nextCycle(1486); checkResult(3123, -2648);
        nextCycle(1487); checkResult(3119, -2653);
        nextCycle(1488); checkResult(3115, -2658);
        nextCycle(1489); checkResult(3111, -2663);
        nextCycle(1490); checkResult(3107, -2668);
        nextCycle(1491); checkResult(3103, -2672);
        nextCycle(1492); checkResult(3099, -2677);
        nextCycle(1493); checkResult(3095, -2682);
        nextCycle(1494); checkResult(3090, -2687);
        nextCycle(1495); checkResult(3086, -2691);
        nextCycle(1496); checkResult(3082, -2696);
        nextCycle(1497); checkResult(3078, -2701);
        nextCycle(1498); checkResult(3074, -2706);
        nextCycle(1499); checkResult(3070, -2710);
        nextCycle(1500); checkResult(3066, -2715);
        nextCycle(1501); checkResult(3061, -2720);
        nextCycle(1502); checkResult(3057, -2724);
        nextCycle(1503); checkResult(3053, -2729);
        nextCycle(1504); checkResult(3049, -2734);
        nextCycle(1505); checkResult(3045, -2738);
        nextCycle(1506); checkResult(3041, -2743);
        nextCycle(1507); checkResult(3036, -2748);
        nextCycle(1508); checkResult(3032, -2752);
        nextCycle(1509); checkResult(3028, -2757);
        nextCycle(1510); checkResult(3024, -2762);
        nextCycle(1511); checkResult(3019, -2766);
        nextCycle(1512); checkResult(3015, -2771);
        nextCycle(1513); checkResult(3011, -2776);
        nextCycle(1514); checkResult(3007, -2780);
        nextCycle(1515); checkResult(3002, -2785);
        nextCycle(1516); checkResult(2998, -2789);
        nextCycle(1517); checkResult(2994, -2794);
        nextCycle(1518); checkResult(2990, -2799);
        nextCycle(1519); checkResult(2985, -2803);
        nextCycle(1520); checkResult(2981, -2808);
        nextCycle(1521); checkResult(2977, -2812);
        nextCycle(1522); checkResult(2972, -2817);
        nextCycle(1523); checkResult(2968, -2821);
        nextCycle(1524); checkResult(2964, -2826);
        nextCycle(1525); checkResult(2959, -2830);
        nextCycle(1526); checkResult(2955, -2835);
        nextCycle(1527); checkResult(2951, -2840);
        nextCycle(1528); checkResult(2946, -2844);
        nextCycle(1529); checkResult(2942, -2849);
        nextCycle(1530); checkResult(2937, -2853);
        nextCycle(1531); checkResult(2933, -2858);
        nextCycle(1532); checkResult(2929, -2862);
        nextCycle(1533); checkResult(2924, -2867);
        nextCycle(1534); checkResult(2920, -2871);
        nextCycle(1535); checkResult(2916, -2876);
        nextCycle(1536); checkResult(2911, -2880);
        nextCycle(1537); checkResult(2907, -2884);
        nextCycle(1538); checkResult(2902, -2889);
        nextCycle(1539); checkResult(2898, -2893);
        nextCycle(1540); checkResult(2893, -2898);
        nextCycle(1541); checkResult(2889, -2902);
        nextCycle(1542); checkResult(2884, -2907);
        nextCycle(1543); checkResult(2880, -2911);
        nextCycle(1544); checkResult(2876, -2916);
        nextCycle(1545); checkResult(2871, -2920);
        nextCycle(1546); checkResult(2867, -2924);
        nextCycle(1547); checkResult(2862, -2929);
        nextCycle(1548); checkResult(2858, -2933);
        nextCycle(1549); checkResult(2853, -2937);
        nextCycle(1550); checkResult(2849, -2942);
        nextCycle(1551); checkResult(2844, -2946);
        nextCycle(1552); checkResult(2840, -2951);
        nextCycle(1553); checkResult(2835, -2955);
        nextCycle(1554); checkResult(2830, -2959);
        nextCycle(1555); checkResult(2826, -2964);
        nextCycle(1556); checkResult(2821, -2968);
        nextCycle(1557); checkResult(2817, -2972);
        nextCycle(1558); checkResult(2812, -2977);
        nextCycle(1559); checkResult(2808, -2981);
        nextCycle(1560); checkResult(2803, -2985);
        nextCycle(1561); checkResult(2799, -2990);
        nextCycle(1562); checkResult(2794, -2994);
        nextCycle(1563); checkResult(2789, -2998);
        nextCycle(1564); checkResult(2785, -3002);
        nextCycle(1565); checkResult(2780, -3007);
        nextCycle(1566); checkResult(2776, -3011);
        nextCycle(1567); checkResult(2771, -3015);
        nextCycle(1568); checkResult(2766, -3019);
        nextCycle(1569); checkResult(2762, -3024);
        nextCycle(1570); checkResult(2757, -3028);
        nextCycle(1571); checkResult(2752, -3032);
        nextCycle(1572); checkResult(2748, -3036);
        nextCycle(1573); checkResult(2743, -3041);
        nextCycle(1574); checkResult(2738, -3045);
        nextCycle(1575); checkResult(2734, -3049);
        nextCycle(1576); checkResult(2729, -3053);
        nextCycle(1577); checkResult(2724, -3057);
        nextCycle(1578); checkResult(2720, -3061);
        nextCycle(1579); checkResult(2715, -3066);
        nextCycle(1580); checkResult(2710, -3070);
        nextCycle(1581); checkResult(2706, -3074);
        nextCycle(1582); checkResult(2701, -3078);
        nextCycle(1583); checkResult(2696, -3082);
        nextCycle(1584); checkResult(2691, -3086);
        nextCycle(1585); checkResult(2687, -3090);
        nextCycle(1586); checkResult(2682, -3095);
        nextCycle(1587); checkResult(2677, -3099);
        nextCycle(1588); checkResult(2672, -3103);
        nextCycle(1589); checkResult(2668, -3107);
        nextCycle(1590); checkResult(2663, -3111);
        nextCycle(1591); checkResult(2658, -3115);
        nextCycle(1592); checkResult(2653, -3119);
        nextCycle(1593); checkResult(2648, -3123);
        nextCycle(1594); checkResult(2644, -3127);
        nextCycle(1595); checkResult(2639, -3131);
        nextCycle(1596); checkResult(2634, -3135);
        nextCycle(1597); checkResult(2629, -3139);
        nextCycle(1598); checkResult(2624, -3143);
        nextCycle(1599); checkResult(2620, -3147);
        nextCycle(1600); checkResult(2615, -3151);
        nextCycle(1601); checkResult(2610, -3155);
        nextCycle(1602); checkResult(2605, -3159);
        nextCycle(1603); checkResult(2600, -3163);
        nextCycle(1604); checkResult(2595, -3167);
        nextCycle(1605); checkResult(2591, -3171);
        nextCycle(1606); checkResult(2586, -3175);
        nextCycle(1607); checkResult(2581, -3179);
        nextCycle(1608); checkResult(2576, -3183);
        nextCycle(1609); checkResult(2571, -3187);
        nextCycle(1610); checkResult(2566, -3191);
        nextCycle(1611); checkResult(2561, -3195);
        nextCycle(1612); checkResult(2556, -3199);
        nextCycle(1613); checkResult(2551, -3203);
        nextCycle(1614); checkResult(2547, -3207);
        nextCycle(1615); checkResult(2542, -3211);
        nextCycle(1616); checkResult(2537, -3215);
        nextCycle(1617); checkResult(2532, -3219);
        nextCycle(1618); checkResult(2527, -3222);
        nextCycle(1619); checkResult(2522, -3226);
        nextCycle(1620); checkResult(2517, -3230);
        nextCycle(1621); checkResult(2512, -3234);
        nextCycle(1622); checkResult(2507, -3238);
        nextCycle(1623); checkResult(2502, -3242);
        nextCycle(1624); checkResult(2497, -3246);
        nextCycle(1625); checkResult(2492, -3249);
        nextCycle(1626); checkResult(2487, -3253);
        nextCycle(1627); checkResult(2482, -3257);
        nextCycle(1628); checkResult(2477, -3261);
        nextCycle(1629); checkResult(2472, -3265);
        nextCycle(1630); checkResult(2467, -3268);
        nextCycle(1631); checkResult(2462, -3272);
        nextCycle(1632); checkResult(2457, -3276);
        nextCycle(1633); checkResult(2452, -3280);
        nextCycle(1634); checkResult(2447, -3284);
        nextCycle(1635); checkResult(2442, -3287);
        nextCycle(1636); checkResult(2437, -3291);
        nextCycle(1637); checkResult(2432, -3295);
        nextCycle(1638); checkResult(2427, -3298);
        nextCycle(1639); checkResult(2422, -3302);
        nextCycle(1640); checkResult(2417, -3306);
        nextCycle(1641); checkResult(2412, -3310);
        nextCycle(1642); checkResult(2406, -3313);
        nextCycle(1643); checkResult(2401, -3317);
        nextCycle(1644); checkResult(2396, -3321);
        nextCycle(1645); checkResult(2391, -3324);
        nextCycle(1646); checkResult(2386, -3328);
        nextCycle(1647); checkResult(2381, -3332);
        nextCycle(1648); checkResult(2376, -3335);
        nextCycle(1649); checkResult(2371, -3339);
        nextCycle(1650); checkResult(2366, -3343);
        nextCycle(1651); checkResult(2361, -3346);
        nextCycle(1652); checkResult(2355, -3350);
        nextCycle(1653); checkResult(2350, -3353);
        nextCycle(1654); checkResult(2345, -3357);
        nextCycle(1655); checkResult(2340, -3361);
        nextCycle(1656); checkResult(2335, -3364);
        nextCycle(1657); checkResult(2330, -3368);
        nextCycle(1658); checkResult(2324, -3371);
        nextCycle(1659); checkResult(2319, -3375);
        nextCycle(1660); checkResult(2314, -3378);
        nextCycle(1661); checkResult(2309, -3382);
        nextCycle(1662); checkResult(2304, -3386);
        nextCycle(1663); checkResult(2299, -3389);
        nextCycle(1664); checkResult(2293, -3393);
        nextCycle(1665); checkResult(2288, -3396);
        nextCycle(1666); checkResult(2283, -3400);
        nextCycle(1667); checkResult(2278, -3403);
        nextCycle(1668); checkResult(2272, -3407);
        nextCycle(1669); checkResult(2267, -3410);
        nextCycle(1670); checkResult(2262, -3414);
        nextCycle(1671); checkResult(2257, -3417);
        nextCycle(1672); checkResult(2252, -3420);
        nextCycle(1673); checkResult(2246, -3424);
        nextCycle(1674); checkResult(2241, -3427);
        nextCycle(1675); checkResult(2236, -3431);
        nextCycle(1676); checkResult(2230, -3434);
        nextCycle(1677); checkResult(2225, -3438);
        nextCycle(1678); checkResult(2220, -3441);
        nextCycle(1679); checkResult(2215, -3444);
        nextCycle(1680); checkResult(2209, -3448);
        nextCycle(1681); checkResult(2204, -3451);
        nextCycle(1682); checkResult(2199, -3455);
        nextCycle(1683); checkResult(2193, -3458);
        nextCycle(1684); checkResult(2188, -3461);
        nextCycle(1685); checkResult(2183, -3465);
        nextCycle(1686); checkResult(2178, -3468);
        nextCycle(1687); checkResult(2172, -3471);
        nextCycle(1688); checkResult(2167, -3475);
        nextCycle(1689); checkResult(2162, -3478);
        nextCycle(1690); checkResult(2156, -3481);
        nextCycle(1691); checkResult(2151, -3485);
        nextCycle(1692); checkResult(2146, -3488);
        nextCycle(1693); checkResult(2140, -3491);
        nextCycle(1694); checkResult(2135, -3495);
        nextCycle(1695); checkResult(2129, -3498);
        nextCycle(1696); checkResult(2124, -3501);
        nextCycle(1697); checkResult(2119, -3504);
        nextCycle(1698); checkResult(2113, -3508);
        nextCycle(1699); checkResult(2108, -3511);
        nextCycle(1700); checkResult(2103, -3514);
        nextCycle(1701); checkResult(2097, -3517);
        nextCycle(1702); checkResult(2092, -3520);
        nextCycle(1703); checkResult(2086, -3524);
        nextCycle(1704); checkResult(2081, -3527);
        nextCycle(1705); checkResult(2076, -3530);
        nextCycle(1706); checkResult(2070, -3533);
        nextCycle(1707); checkResult(2065, -3536);
        nextCycle(1708); checkResult(2059, -3540);
        nextCycle(1709); checkResult(2054, -3543);
        nextCycle(1710); checkResult(2048, -3546);
        nextCycle(1711); checkResult(2043, -3549);
        nextCycle(1712); checkResult(2038, -3552);
        nextCycle(1713); checkResult(2032, -3555);
        nextCycle(1714); checkResult(2027, -3558);
        nextCycle(1715); checkResult(2021, -3561);
        nextCycle(1716); checkResult(2016, -3565);
        nextCycle(1717); checkResult(2010, -3568);
        nextCycle(1718); checkResult(2005, -3571);
        nextCycle(1719); checkResult(1999, -3574);
        nextCycle(1720); checkResult(1994, -3577);
        nextCycle(1721); checkResult(1988, -3580);
        nextCycle(1722); checkResult(1983, -3583);
        nextCycle(1723); checkResult(1977, -3586);
        nextCycle(1724); checkResult(1972, -3589);
        nextCycle(1725); checkResult(1966, -3592);
        nextCycle(1726); checkResult(1961, -3595);
        nextCycle(1727); checkResult(1955, -3598);
        nextCycle(1728); checkResult(1950, -3601);
        nextCycle(1729); checkResult(1944, -3604);
        nextCycle(1730); checkResult(1939, -3607);
        nextCycle(1731); checkResult(1933, -3610);
        nextCycle(1732); checkResult(1928, -3613);
        nextCycle(1733); checkResult(1922, -3616);
        nextCycle(1734); checkResult(1917, -3619);
        nextCycle(1735); checkResult(1911, -3622);
        nextCycle(1736); checkResult(1905, -3625);
        nextCycle(1737); checkResult(1900, -3628);
        nextCycle(1738); checkResult(1894, -3631);
        nextCycle(1739); checkResult(1889, -3633);
        nextCycle(1740); checkResult(1883, -3636);
        nextCycle(1741); checkResult(1878, -3639);
        nextCycle(1742); checkResult(1872, -3642);
        nextCycle(1743); checkResult(1866, -3645);
        nextCycle(1744); checkResult(1861, -3648);
        nextCycle(1745); checkResult(1855, -3651);
        nextCycle(1746); checkResult(1850, -3654);
        nextCycle(1747); checkResult(1844, -3656);
        nextCycle(1748); checkResult(1838, -3659);
        nextCycle(1749); checkResult(1833, -3662);
        nextCycle(1750); checkResult(1827, -3665);
        nextCycle(1751); checkResult(1821, -3668);
        nextCycle(1752); checkResult(1816, -3670);
        nextCycle(1753); checkResult(1810, -3673);
        nextCycle(1754); checkResult(1805, -3676);
        nextCycle(1755); checkResult(1799, -3679);
        nextCycle(1756); checkResult(1793, -3681);
        nextCycle(1757); checkResult(1788, -3684);
        nextCycle(1758); checkResult(1782, -3687);
        nextCycle(1759); checkResult(1776, -3690);
        nextCycle(1760); checkResult(1771, -3692);
        nextCycle(1761); checkResult(1765, -3695);
        nextCycle(1762); checkResult(1759, -3698);
        nextCycle(1763); checkResult(1754, -3700);
        nextCycle(1764); checkResult(1748, -3703);
        nextCycle(1765); checkResult(1742, -3706);
        nextCycle(1766); checkResult(1737, -3709);
        nextCycle(1767); checkResult(1731, -3711);
        nextCycle(1768); checkResult(1725, -3714);
        nextCycle(1769); checkResult(1720, -3716);
        nextCycle(1770); checkResult(1714, -3719);
        nextCycle(1771); checkResult(1708, -3722);
        nextCycle(1772); checkResult(1702, -3724);
        nextCycle(1773); checkResult(1697, -3727);
        nextCycle(1774); checkResult(1691, -3730);
        nextCycle(1775); checkResult(1685, -3732);
        nextCycle(1776); checkResult(1680, -3735);
        nextCycle(1777); checkResult(1674, -3737);
        nextCycle(1778); checkResult(1668, -3740);
        nextCycle(1779); checkResult(1662, -3742);
        nextCycle(1780); checkResult(1657, -3745);
        nextCycle(1781); checkResult(1651, -3747);
        nextCycle(1782); checkResult(1645, -3750);
        nextCycle(1783); checkResult(1639, -3753);
        nextCycle(1784); checkResult(1634, -3755);
        nextCycle(1785); checkResult(1628, -3758);
        nextCycle(1786); checkResult(1622, -3760);
        nextCycle(1787); checkResult(1616, -3763);
        nextCycle(1788); checkResult(1611, -3765);
        nextCycle(1789); checkResult(1605, -3767);
        nextCycle(1790); checkResult(1599, -3770);
        nextCycle(1791); checkResult(1593, -3772);
        nextCycle(1792); checkResult(1587, -3775);
        nextCycle(1793); checkResult(1582, -3777);
        nextCycle(1794); checkResult(1576, -3780);
        nextCycle(1795); checkResult(1570, -3782);
        nextCycle(1796); checkResult(1564, -3784);
        nextCycle(1797); checkResult(1558, -3787);
        nextCycle(1798); checkResult(1553, -3789);
        nextCycle(1799); checkResult(1547, -3792);
        nextCycle(1800); checkResult(1541, -3794);
        nextCycle(1801); checkResult(1535, -3796);
        nextCycle(1802); checkResult(1529, -3799);
        nextCycle(1803); checkResult(1523, -3801);
        nextCycle(1804); checkResult(1518, -3803);
        nextCycle(1805); checkResult(1512, -3806);
        nextCycle(1806); checkResult(1506, -3808);
        nextCycle(1807); checkResult(1500, -3810);
        nextCycle(1808); checkResult(1494, -3813);
        nextCycle(1809); checkResult(1488, -3815);
        nextCycle(1810); checkResult(1483, -3817);
        nextCycle(1811); checkResult(1477, -3819);
        nextCycle(1812); checkResult(1471, -3822);
        nextCycle(1813); checkResult(1465, -3824);
        nextCycle(1814); checkResult(1459, -3826);
        nextCycle(1815); checkResult(1453, -3828);
        nextCycle(1816); checkResult(1447, -3831);
        nextCycle(1817); checkResult(1441, -3833);
        nextCycle(1818); checkResult(1436, -3835);
        nextCycle(1819); checkResult(1430, -3837);
        nextCycle(1820); checkResult(1424, -3839);
        nextCycle(1821); checkResult(1418, -3842);
        nextCycle(1822); checkResult(1412, -3844);
        nextCycle(1823); checkResult(1406, -3846);
        nextCycle(1824); checkResult(1400, -3848);
        nextCycle(1825); checkResult(1394, -3850);
        nextCycle(1826); checkResult(1388, -3852);
        nextCycle(1827); checkResult(1383, -3855);
        nextCycle(1828); checkResult(1377, -3857);
        nextCycle(1829); checkResult(1371, -3859);
        nextCycle(1830); checkResult(1365, -3861);
        nextCycle(1831); checkResult(1359, -3863);
        nextCycle(1832); checkResult(1353, -3865);
        nextCycle(1833); checkResult(1347, -3867);
        nextCycle(1834); checkResult(1341, -3869);
        nextCycle(1835); checkResult(1335, -3871);
        nextCycle(1836); checkResult(1329, -3873);
        nextCycle(1837); checkResult(1323, -3875);
        nextCycle(1838); checkResult(1317, -3877);
        nextCycle(1839); checkResult(1311, -3879);
        nextCycle(1840); checkResult(1305, -3881);
        nextCycle(1841); checkResult(1299, -3883);
        nextCycle(1842); checkResult(1293, -3885);
        nextCycle(1843); checkResult(1288, -3887);
        nextCycle(1844); checkResult(1282, -3889);
        nextCycle(1845); checkResult(1276, -3891);
        nextCycle(1846); checkResult(1270, -3893);
        nextCycle(1847); checkResult(1264, -3895);
        nextCycle(1848); checkResult(1258, -3897);
        nextCycle(1849); checkResult(1252, -3899);
        nextCycle(1850); checkResult(1246, -3901);
        nextCycle(1851); checkResult(1240, -3903);
        nextCycle(1852); checkResult(1234, -3905);
        nextCycle(1853); checkResult(1228, -3907);
        nextCycle(1854); checkResult(1222, -3909);
        nextCycle(1855); checkResult(1216, -3910);
        nextCycle(1856); checkResult(1210, -3912);
        nextCycle(1857); checkResult(1204, -3914);
        nextCycle(1858); checkResult(1198, -3916);
        nextCycle(1859); checkResult(1192, -3918);
        nextCycle(1860); checkResult(1186, -3920);
        nextCycle(1861); checkResult(1180, -3921);
        nextCycle(1862); checkResult(1174, -3923);
        nextCycle(1863); checkResult(1168, -3925);
        nextCycle(1864); checkResult(1162, -3927);
        nextCycle(1865); checkResult(1156, -3929);
        nextCycle(1866); checkResult(1150, -3930);
        nextCycle(1867); checkResult(1144, -3932);
        nextCycle(1868); checkResult(1138, -3934);
        nextCycle(1869); checkResult(1131, -3936);
        nextCycle(1870); checkResult(1125, -3937);
        nextCycle(1871); checkResult(1119, -3939);
        nextCycle(1872); checkResult(1113, -3941);
        nextCycle(1873); checkResult(1107, -3942);
        nextCycle(1874); checkResult(1101, -3944);
        nextCycle(1875); checkResult(1095, -3946);
        nextCycle(1876); checkResult(1089, -3947);
        nextCycle(1877); checkResult(1083, -3949);
        nextCycle(1878); checkResult(1077, -3951);
        nextCycle(1879); checkResult(1071, -3952);
        nextCycle(1880); checkResult(1065, -3954);
        nextCycle(1881); checkResult(1059, -3956);
        nextCycle(1882); checkResult(1053, -3957);
        nextCycle(1883); checkResult(1047, -3959);
        nextCycle(1884); checkResult(1041, -3961);
        nextCycle(1885); checkResult(1035, -3962);
        nextCycle(1886); checkResult(1028, -3964);
        nextCycle(1887); checkResult(1022, -3965);
        nextCycle(1888); checkResult(1016, -3967);
        nextCycle(1889); checkResult(1010, -3968);
        nextCycle(1890); checkResult(1004, -3970);
        nextCycle(1891); checkResult(998, -3972);
        nextCycle(1892); checkResult(992, -3973);
        nextCycle(1893); checkResult(986, -3975);
        nextCycle(1894); checkResult(980, -3976);
        nextCycle(1895); checkResult(974, -3978);
        nextCycle(1896); checkResult(968, -3979);
        nextCycle(1897); checkResult(961, -3981);
        nextCycle(1898); checkResult(955, -3982);
        nextCycle(1899); checkResult(949, -3983);
        nextCycle(1900); checkResult(943, -3985);
        nextCycle(1901); checkResult(937, -3986);
        nextCycle(1902); checkResult(931, -3988);
        nextCycle(1903); checkResult(925, -3989);
        nextCycle(1904); checkResult(919, -3991);
        nextCycle(1905); checkResult(913, -3992);
        nextCycle(1906); checkResult(906, -3993);
        nextCycle(1907); checkResult(900, -3995);
        nextCycle(1908); checkResult(894, -3996);
        nextCycle(1909); checkResult(888, -3998);
        nextCycle(1910); checkResult(882, -3999);
        nextCycle(1911); checkResult(876, -4000);
        nextCycle(1912); checkResult(870, -4002);
        nextCycle(1913); checkResult(863, -4003);
        nextCycle(1914); checkResult(857, -4004);
        nextCycle(1915); checkResult(851, -4006);
        nextCycle(1916); checkResult(845, -4007);
        nextCycle(1917); checkResult(839, -4008);
        nextCycle(1918); checkResult(833, -4009);
        nextCycle(1919); checkResult(827, -4011);
        nextCycle(1920); checkResult(820, -4012);
        nextCycle(1921); checkResult(814, -4013);
        nextCycle(1922); checkResult(808, -4014);
        nextCycle(1923); checkResult(802, -4016);
        nextCycle(1924); checkResult(796, -4017);
        nextCycle(1925); checkResult(790, -4018);
        nextCycle(1926); checkResult(783, -4019);
        nextCycle(1927); checkResult(777, -4021);
        nextCycle(1928); checkResult(771, -4022);
        nextCycle(1929); checkResult(765, -4023);
        nextCycle(1930); checkResult(759, -4024);
        nextCycle(1931); checkResult(753, -4025);
        nextCycle(1932); checkResult(746, -4026);
        nextCycle(1933); checkResult(740, -4028);
        nextCycle(1934); checkResult(734, -4029);
        nextCycle(1935); checkResult(728, -4030);
        nextCycle(1936); checkResult(722, -4031);
        nextCycle(1937); checkResult(716, -4032);
        nextCycle(1938); checkResult(709, -4033);
        nextCycle(1939); checkResult(703, -4034);
        nextCycle(1940); checkResult(697, -4035);
        nextCycle(1941); checkResult(691, -4036);
        nextCycle(1942); checkResult(685, -4037);
        nextCycle(1943); checkResult(678, -4038);
        nextCycle(1944); checkResult(672, -4039);
        nextCycle(1945); checkResult(666, -4040);
        nextCycle(1946); checkResult(660, -4041);
        nextCycle(1947); checkResult(654, -4042);
        nextCycle(1948); checkResult(647, -4043);
        nextCycle(1949); checkResult(641, -4044);
        nextCycle(1950); checkResult(635, -4045);
        nextCycle(1951); checkResult(629, -4046);
        nextCycle(1952); checkResult(623, -4047);
        nextCycle(1953); checkResult(616, -4048);
        nextCycle(1954); checkResult(610, -4049);
        nextCycle(1955); checkResult(604, -4050);
        nextCycle(1956); checkResult(598, -4051);
        nextCycle(1957); checkResult(592, -4052);
        nextCycle(1958); checkResult(585, -4053);
        nextCycle(1959); checkResult(579, -4054);
        nextCycle(1960); checkResult(573, -4055);
        nextCycle(1961); checkResult(567, -4056);
        nextCycle(1962); checkResult(560, -4056);
        nextCycle(1963); checkResult(554, -4057);
        nextCycle(1964); checkResult(548, -4058);
        nextCycle(1965); checkResult(542, -4059);
        nextCycle(1966); checkResult(536, -4060);
        nextCycle(1967); checkResult(529, -4061);
        nextCycle(1968); checkResult(523, -4061);
        nextCycle(1969); checkResult(517, -4062);
        nextCycle(1970); checkResult(511, -4063);
        nextCycle(1971); checkResult(504, -4064);
        nextCycle(1972); checkResult(498, -4065);
        nextCycle(1973); checkResult(492, -4065);
        nextCycle(1974); checkResult(486, -4066);
        nextCycle(1975); checkResult(479, -4067);
        nextCycle(1976); checkResult(473, -4068);
        nextCycle(1977); checkResult(467, -4068);
        nextCycle(1978); checkResult(461, -4069);
        nextCycle(1979); checkResult(454, -4070);
        nextCycle(1980); checkResult(448, -4070);
        nextCycle(1981); checkResult(442, -4071);
        nextCycle(1982); checkResult(436, -4072);
        nextCycle(1983); checkResult(430, -4072);
        nextCycle(1984); checkResult(423, -4073);
        nextCycle(1985); checkResult(417, -4074);
        nextCycle(1986); checkResult(411, -4074);
        nextCycle(1987); checkResult(405, -4075);
        nextCycle(1988); checkResult(398, -4076);
        nextCycle(1989); checkResult(392, -4076);
        nextCycle(1990); checkResult(386, -4077);
        nextCycle(1991); checkResult(379, -4077);
        nextCycle(1992); checkResult(373, -4078);
        nextCycle(1993); checkResult(367, -4079);
        nextCycle(1994); checkResult(361, -4079);
        nextCycle(1995); checkResult(354, -4080);
        nextCycle(1996); checkResult(348, -4080);
        nextCycle(1997); checkResult(342, -4081);
        nextCycle(1998); checkResult(336, -4081);
        nextCycle(1999); checkResult(329, -4082);
        nextCycle(2000); checkResult(323, -4082);
        nextCycle(2001); checkResult(317, -4083);
        nextCycle(2002); checkResult(311, -4083);
        nextCycle(2003); checkResult(304, -4084);
        nextCycle(2004); checkResult(298, -4084);
        nextCycle(2005); checkResult(292, -4085);
        nextCycle(2006); checkResult(286, -4085);
        nextCycle(2007); checkResult(279, -4085);
        nextCycle(2008); checkResult(273, -4086);
        nextCycle(2009); checkResult(267, -4086);
        nextCycle(2010); checkResult(261, -4087);
        nextCycle(2011); checkResult(254, -4087);
        nextCycle(2012); checkResult(248, -4087);
        nextCycle(2013); checkResult(242, -4088);
        nextCycle(2014); checkResult(235, -4088);
        nextCycle(2015); checkResult(229, -4089);
        nextCycle(2016); checkResult(223, -4089);
        nextCycle(2017); checkResult(217, -4089);
        nextCycle(2018); checkResult(210, -4090);
        nextCycle(2019); checkResult(204, -4090);
        nextCycle(2020); checkResult(198, -4090);
        nextCycle(2021); checkResult(192, -4091);
        nextCycle(2022); checkResult(185, -4091);
        nextCycle(2023); checkResult(179, -4091);
        nextCycle(2024); checkResult(173, -4091);
        nextCycle(2025); checkResult(166, -4092);
        nextCycle(2026); checkResult(160, -4092);
        nextCycle(2027); checkResult(154, -4092);
        nextCycle(2028); checkResult(148, -4092);
        nextCycle(2029); checkResult(141, -4093);
        nextCycle(2030); checkResult(135, -4093);
        nextCycle(2031); checkResult(129, -4093);
        nextCycle(2032); checkResult(122, -4093);
        nextCycle(2033); checkResult(116, -4093);
        nextCycle(2034); checkResult(110, -4094);
        nextCycle(2035); checkResult(104, -4094);
        nextCycle(2036); checkResult(97, -4094);
        nextCycle(2037); checkResult(91, -4094);
        nextCycle(2038); checkResult(85, -4094);
        nextCycle(2039); checkResult(79, -4094);
        nextCycle(2040); checkResult(72, -4094);
        nextCycle(2041); checkResult(66, -4094);
        nextCycle(2042); checkResult(60, -4095);
        nextCycle(2043); checkResult(53, -4095);
        nextCycle(2044); checkResult(47, -4095);
        nextCycle(2045); checkResult(41, -4095);
        nextCycle(2046); checkResult(35, -4095);
        nextCycle(2047); checkResult(28, -4095);
        nextCycle(2048); checkResult(22, -4095);
        nextCycle(2049); checkResult(16, -4095);
        nextCycle(2050); checkResult(9, -4095);
        nextCycle(2051); checkResult(3, -4095);
        nextCycle(2052); checkResult(-3, -4095);
        nextCycle(2053); checkResult(-9, -4095);
        nextCycle(2054); checkResult(-16, -4095);
        nextCycle(2055); checkResult(-22, -4095);
        nextCycle(2056); checkResult(-28, -4095);
        nextCycle(2057); checkResult(-35, -4095);
        nextCycle(2058); checkResult(-41, -4095);
        nextCycle(2059); checkResult(-47, -4095);
        nextCycle(2060); checkResult(-53, -4095);
        nextCycle(2061); checkResult(-60, -4095);
        nextCycle(2062); checkResult(-66, -4094);
        nextCycle(2063); checkResult(-72, -4094);
        nextCycle(2064); checkResult(-79, -4094);
        nextCycle(2065); checkResult(-85, -4094);
        nextCycle(2066); checkResult(-91, -4094);
        nextCycle(2067); checkResult(-97, -4094);
        nextCycle(2068); checkResult(-104, -4094);
        nextCycle(2069); checkResult(-110, -4094);
        nextCycle(2070); checkResult(-116, -4093);
        nextCycle(2071); checkResult(-122, -4093);
        nextCycle(2072); checkResult(-129, -4093);
        nextCycle(2073); checkResult(-135, -4093);
        nextCycle(2074); checkResult(-141, -4093);
        nextCycle(2075); checkResult(-148, -4092);
        nextCycle(2076); checkResult(-154, -4092);
        nextCycle(2077); checkResult(-160, -4092);
        nextCycle(2078); checkResult(-166, -4092);
        nextCycle(2079); checkResult(-173, -4091);
        nextCycle(2080); checkResult(-179, -4091);
        nextCycle(2081); checkResult(-185, -4091);
        nextCycle(2082); checkResult(-192, -4091);
        nextCycle(2083); checkResult(-198, -4090);
        nextCycle(2084); checkResult(-204, -4090);
        nextCycle(2085); checkResult(-210, -4090);
        nextCycle(2086); checkResult(-217, -4089);
        nextCycle(2087); checkResult(-223, -4089);
        nextCycle(2088); checkResult(-229, -4089);
        nextCycle(2089); checkResult(-235, -4088);
        nextCycle(2090); checkResult(-242, -4088);
        nextCycle(2091); checkResult(-248, -4087);
        nextCycle(2092); checkResult(-254, -4087);
        nextCycle(2093); checkResult(-261, -4087);
        nextCycle(2094); checkResult(-267, -4086);
        nextCycle(2095); checkResult(-273, -4086);
        nextCycle(2096); checkResult(-279, -4085);
        nextCycle(2097); checkResult(-286, -4085);
        nextCycle(2098); checkResult(-292, -4085);
        nextCycle(2099); checkResult(-298, -4084);
        nextCycle(2100); checkResult(-304, -4084);
        nextCycle(2101); checkResult(-311, -4083);
        nextCycle(2102); checkResult(-317, -4083);
        nextCycle(2103); checkResult(-323, -4082);
        nextCycle(2104); checkResult(-329, -4082);
        nextCycle(2105); checkResult(-336, -4081);
        nextCycle(2106); checkResult(-342, -4081);
        nextCycle(2107); checkResult(-348, -4080);
        nextCycle(2108); checkResult(-354, -4080);
        nextCycle(2109); checkResult(-361, -4079);
        nextCycle(2110); checkResult(-367, -4079);
        nextCycle(2111); checkResult(-373, -4078);
        nextCycle(2112); checkResult(-379, -4077);
        nextCycle(2113); checkResult(-386, -4077);
        nextCycle(2114); checkResult(-392, -4076);
        nextCycle(2115); checkResult(-398, -4076);
        nextCycle(2116); checkResult(-405, -4075);
        nextCycle(2117); checkResult(-411, -4074);
        nextCycle(2118); checkResult(-417, -4074);
        nextCycle(2119); checkResult(-423, -4073);
        nextCycle(2120); checkResult(-430, -4072);
        nextCycle(2121); checkResult(-436, -4072);
        nextCycle(2122); checkResult(-442, -4071);
        nextCycle(2123); checkResult(-448, -4070);
        nextCycle(2124); checkResult(-454, -4070);
        nextCycle(2125); checkResult(-461, -4069);
        nextCycle(2126); checkResult(-467, -4068);
        nextCycle(2127); checkResult(-473, -4068);
        nextCycle(2128); checkResult(-479, -4067);
        nextCycle(2129); checkResult(-486, -4066);
        nextCycle(2130); checkResult(-492, -4065);
        nextCycle(2131); checkResult(-498, -4065);
        nextCycle(2132); checkResult(-504, -4064);
        nextCycle(2133); checkResult(-511, -4063);
        nextCycle(2134); checkResult(-517, -4062);
        nextCycle(2135); checkResult(-523, -4061);
        nextCycle(2136); checkResult(-529, -4061);
        nextCycle(2137); checkResult(-536, -4060);
        nextCycle(2138); checkResult(-542, -4059);
        nextCycle(2139); checkResult(-548, -4058);
        nextCycle(2140); checkResult(-554, -4057);
        nextCycle(2141); checkResult(-560, -4056);
        nextCycle(2142); checkResult(-567, -4056);
        nextCycle(2143); checkResult(-573, -4055);
        nextCycle(2144); checkResult(-579, -4054);
        nextCycle(2145); checkResult(-585, -4053);
        nextCycle(2146); checkResult(-592, -4052);
        nextCycle(2147); checkResult(-598, -4051);
        nextCycle(2148); checkResult(-604, -4050);
        nextCycle(2149); checkResult(-610, -4049);
        nextCycle(2150); checkResult(-616, -4048);
        nextCycle(2151); checkResult(-623, -4047);
        nextCycle(2152); checkResult(-629, -4046);
        nextCycle(2153); checkResult(-635, -4045);
        nextCycle(2154); checkResult(-641, -4044);
        nextCycle(2155); checkResult(-647, -4043);
        nextCycle(2156); checkResult(-654, -4042);
        nextCycle(2157); checkResult(-660, -4041);
        nextCycle(2158); checkResult(-666, -4040);
        nextCycle(2159); checkResult(-672, -4039);
        nextCycle(2160); checkResult(-678, -4038);
        nextCycle(2161); checkResult(-685, -4037);
        nextCycle(2162); checkResult(-691, -4036);
        nextCycle(2163); checkResult(-697, -4035);
        nextCycle(2164); checkResult(-703, -4034);
        nextCycle(2165); checkResult(-709, -4033);
        nextCycle(2166); checkResult(-716, -4032);
        nextCycle(2167); checkResult(-722, -4031);
        nextCycle(2168); checkResult(-728, -4030);
        nextCycle(2169); checkResult(-734, -4029);
        nextCycle(2170); checkResult(-740, -4028);
        nextCycle(2171); checkResult(-746, -4026);
        nextCycle(2172); checkResult(-753, -4025);
        nextCycle(2173); checkResult(-759, -4024);
        nextCycle(2174); checkResult(-765, -4023);
        nextCycle(2175); checkResult(-771, -4022);
        nextCycle(2176); checkResult(-777, -4021);
        nextCycle(2177); checkResult(-783, -4019);
        nextCycle(2178); checkResult(-790, -4018);
        nextCycle(2179); checkResult(-796, -4017);
        nextCycle(2180); checkResult(-802, -4016);
        nextCycle(2181); checkResult(-808, -4014);
        nextCycle(2182); checkResult(-814, -4013);
        nextCycle(2183); checkResult(-820, -4012);
        nextCycle(2184); checkResult(-827, -4011);
        nextCycle(2185); checkResult(-833, -4009);
        nextCycle(2186); checkResult(-839, -4008);
        nextCycle(2187); checkResult(-845, -4007);
        nextCycle(2188); checkResult(-851, -4006);
        nextCycle(2189); checkResult(-857, -4004);
        nextCycle(2190); checkResult(-863, -4003);
        nextCycle(2191); checkResult(-870, -4002);
        nextCycle(2192); checkResult(-876, -4000);
        nextCycle(2193); checkResult(-882, -3999);
        nextCycle(2194); checkResult(-888, -3998);
        nextCycle(2195); checkResult(-894, -3996);
        nextCycle(2196); checkResult(-900, -3995);
        nextCycle(2197); checkResult(-906, -3993);
        nextCycle(2198); checkResult(-913, -3992);
        nextCycle(2199); checkResult(-919, -3991);
        nextCycle(2200); checkResult(-925, -3989);
        nextCycle(2201); checkResult(-931, -3988);
        nextCycle(2202); checkResult(-937, -3986);
        nextCycle(2203); checkResult(-943, -3985);
        nextCycle(2204); checkResult(-949, -3983);
        nextCycle(2205); checkResult(-955, -3982);
        nextCycle(2206); checkResult(-961, -3981);
        nextCycle(2207); checkResult(-968, -3979);
        nextCycle(2208); checkResult(-974, -3978);
        nextCycle(2209); checkResult(-980, -3976);
        nextCycle(2210); checkResult(-986, -3975);
        nextCycle(2211); checkResult(-992, -3973);
        nextCycle(2212); checkResult(-998, -3972);
        nextCycle(2213); checkResult(-1004, -3970);
        nextCycle(2214); checkResult(-1010, -3968);
        nextCycle(2215); checkResult(-1016, -3967);
        nextCycle(2216); checkResult(-1022, -3965);
        nextCycle(2217); checkResult(-1028, -3964);
        nextCycle(2218); checkResult(-1035, -3962);
        nextCycle(2219); checkResult(-1041, -3961);
        nextCycle(2220); checkResult(-1047, -3959);
        nextCycle(2221); checkResult(-1053, -3957);
        nextCycle(2222); checkResult(-1059, -3956);
        nextCycle(2223); checkResult(-1065, -3954);
        nextCycle(2224); checkResult(-1071, -3952);
        nextCycle(2225); checkResult(-1077, -3951);
        nextCycle(2226); checkResult(-1083, -3949);
        nextCycle(2227); checkResult(-1089, -3947);
        nextCycle(2228); checkResult(-1095, -3946);
        nextCycle(2229); checkResult(-1101, -3944);
        nextCycle(2230); checkResult(-1107, -3942);
        nextCycle(2231); checkResult(-1113, -3941);
        nextCycle(2232); checkResult(-1119, -3939);
        nextCycle(2233); checkResult(-1125, -3937);
        nextCycle(2234); checkResult(-1131, -3936);
        nextCycle(2235); checkResult(-1138, -3934);
        nextCycle(2236); checkResult(-1144, -3932);
        nextCycle(2237); checkResult(-1150, -3930);
        nextCycle(2238); checkResult(-1156, -3929);
        nextCycle(2239); checkResult(-1162, -3927);
        nextCycle(2240); checkResult(-1168, -3925);
        nextCycle(2241); checkResult(-1174, -3923);
        nextCycle(2242); checkResult(-1180, -3921);
        nextCycle(2243); checkResult(-1186, -3920);
        nextCycle(2244); checkResult(-1192, -3918);
        nextCycle(2245); checkResult(-1198, -3916);
        nextCycle(2246); checkResult(-1204, -3914);
        nextCycle(2247); checkResult(-1210, -3912);
        nextCycle(2248); checkResult(-1216, -3910);
        nextCycle(2249); checkResult(-1222, -3909);
        nextCycle(2250); checkResult(-1228, -3907);
        nextCycle(2251); checkResult(-1234, -3905);
        nextCycle(2252); checkResult(-1240, -3903);
        nextCycle(2253); checkResult(-1246, -3901);
        nextCycle(2254); checkResult(-1252, -3899);
        nextCycle(2255); checkResult(-1258, -3897);
        nextCycle(2256); checkResult(-1264, -3895);
        nextCycle(2257); checkResult(-1270, -3893);
        nextCycle(2258); checkResult(-1276, -3891);
        nextCycle(2259); checkResult(-1282, -3889);
        nextCycle(2260); checkResult(-1288, -3887);
        nextCycle(2261); checkResult(-1293, -3885);
        nextCycle(2262); checkResult(-1299, -3883);
        nextCycle(2263); checkResult(-1305, -3881);
        nextCycle(2264); checkResult(-1311, -3879);
        nextCycle(2265); checkResult(-1317, -3877);
        nextCycle(2266); checkResult(-1323, -3875);
        nextCycle(2267); checkResult(-1329, -3873);
        nextCycle(2268); checkResult(-1335, -3871);
        nextCycle(2269); checkResult(-1341, -3869);
        nextCycle(2270); checkResult(-1347, -3867);
        nextCycle(2271); checkResult(-1353, -3865);
        nextCycle(2272); checkResult(-1359, -3863);
        nextCycle(2273); checkResult(-1365, -3861);
        nextCycle(2274); checkResult(-1371, -3859);
        nextCycle(2275); checkResult(-1377, -3857);
        nextCycle(2276); checkResult(-1383, -3855);
        nextCycle(2277); checkResult(-1388, -3852);
        nextCycle(2278); checkResult(-1394, -3850);
        nextCycle(2279); checkResult(-1400, -3848);
        nextCycle(2280); checkResult(-1406, -3846);
        nextCycle(2281); checkResult(-1412, -3844);
        nextCycle(2282); checkResult(-1418, -3842);
        nextCycle(2283); checkResult(-1424, -3839);
        nextCycle(2284); checkResult(-1430, -3837);
        nextCycle(2285); checkResult(-1436, -3835);
        nextCycle(2286); checkResult(-1441, -3833);
        nextCycle(2287); checkResult(-1447, -3831);
        nextCycle(2288); checkResult(-1453, -3828);
        nextCycle(2289); checkResult(-1459, -3826);
        nextCycle(2290); checkResult(-1465, -3824);
        nextCycle(2291); checkResult(-1471, -3822);
        nextCycle(2292); checkResult(-1477, -3819);
        nextCycle(2293); checkResult(-1483, -3817);
        nextCycle(2294); checkResult(-1488, -3815);
        nextCycle(2295); checkResult(-1494, -3813);
        nextCycle(2296); checkResult(-1500, -3810);
        nextCycle(2297); checkResult(-1506, -3808);
        nextCycle(2298); checkResult(-1512, -3806);
        nextCycle(2299); checkResult(-1518, -3803);
        nextCycle(2300); checkResult(-1523, -3801);
        nextCycle(2301); checkResult(-1529, -3799);
        nextCycle(2302); checkResult(-1535, -3796);
        nextCycle(2303); checkResult(-1541, -3794);
        nextCycle(2304); checkResult(-1547, -3792);
        nextCycle(2305); checkResult(-1553, -3789);
        nextCycle(2306); checkResult(-1558, -3787);
        nextCycle(2307); checkResult(-1564, -3784);
        nextCycle(2308); checkResult(-1570, -3782);
        nextCycle(2309); checkResult(-1576, -3780);
        nextCycle(2310); checkResult(-1582, -3777);
        nextCycle(2311); checkResult(-1587, -3775);
        nextCycle(2312); checkResult(-1593, -3772);
        nextCycle(2313); checkResult(-1599, -3770);
        nextCycle(2314); checkResult(-1605, -3767);
        nextCycle(2315); checkResult(-1611, -3765);
        nextCycle(2316); checkResult(-1616, -3763);
        nextCycle(2317); checkResult(-1622, -3760);
        nextCycle(2318); checkResult(-1628, -3758);
        nextCycle(2319); checkResult(-1634, -3755);
        nextCycle(2320); checkResult(-1639, -3753);
        nextCycle(2321); checkResult(-1645, -3750);
        nextCycle(2322); checkResult(-1651, -3747);
        nextCycle(2323); checkResult(-1657, -3745);
        nextCycle(2324); checkResult(-1662, -3742);
        nextCycle(2325); checkResult(-1668, -3740);
        nextCycle(2326); checkResult(-1674, -3737);
        nextCycle(2327); checkResult(-1680, -3735);
        nextCycle(2328); checkResult(-1685, -3732);
        nextCycle(2329); checkResult(-1691, -3730);
        nextCycle(2330); checkResult(-1697, -3727);
        nextCycle(2331); checkResult(-1702, -3724);
        nextCycle(2332); checkResult(-1708, -3722);
        nextCycle(2333); checkResult(-1714, -3719);
        nextCycle(2334); checkResult(-1720, -3716);
        nextCycle(2335); checkResult(-1725, -3714);
        nextCycle(2336); checkResult(-1731, -3711);
        nextCycle(2337); checkResult(-1737, -3709);
        nextCycle(2338); checkResult(-1742, -3706);
        nextCycle(2339); checkResult(-1748, -3703);
        nextCycle(2340); checkResult(-1754, -3700);
        nextCycle(2341); checkResult(-1759, -3698);
        nextCycle(2342); checkResult(-1765, -3695);
        nextCycle(2343); checkResult(-1771, -3692);
        nextCycle(2344); checkResult(-1776, -3690);
        nextCycle(2345); checkResult(-1782, -3687);
        nextCycle(2346); checkResult(-1788, -3684);
        nextCycle(2347); checkResult(-1793, -3681);
        nextCycle(2348); checkResult(-1799, -3679);
        nextCycle(2349); checkResult(-1805, -3676);
        nextCycle(2350); checkResult(-1810, -3673);
        nextCycle(2351); checkResult(-1816, -3670);
        nextCycle(2352); checkResult(-1821, -3668);
        nextCycle(2353); checkResult(-1827, -3665);
        nextCycle(2354); checkResult(-1833, -3662);
        nextCycle(2355); checkResult(-1838, -3659);
        nextCycle(2356); checkResult(-1844, -3656);
        nextCycle(2357); checkResult(-1850, -3654);
        nextCycle(2358); checkResult(-1855, -3651);
        nextCycle(2359); checkResult(-1861, -3648);
        nextCycle(2360); checkResult(-1866, -3645);
        nextCycle(2361); checkResult(-1872, -3642);
        nextCycle(2362); checkResult(-1878, -3639);
        nextCycle(2363); checkResult(-1883, -3636);
        nextCycle(2364); checkResult(-1889, -3633);
        nextCycle(2365); checkResult(-1894, -3631);
        nextCycle(2366); checkResult(-1900, -3628);
        nextCycle(2367); checkResult(-1905, -3625);
        nextCycle(2368); checkResult(-1911, -3622);
        nextCycle(2369); checkResult(-1917, -3619);
        nextCycle(2370); checkResult(-1922, -3616);
        nextCycle(2371); checkResult(-1928, -3613);
        nextCycle(2372); checkResult(-1933, -3610);
        nextCycle(2373); checkResult(-1939, -3607);
        nextCycle(2374); checkResult(-1944, -3604);
        nextCycle(2375); checkResult(-1950, -3601);
        nextCycle(2376); checkResult(-1955, -3598);
        nextCycle(2377); checkResult(-1961, -3595);
        nextCycle(2378); checkResult(-1966, -3592);
        nextCycle(2379); checkResult(-1972, -3589);
        nextCycle(2380); checkResult(-1977, -3586);
        nextCycle(2381); checkResult(-1983, -3583);
        nextCycle(2382); checkResult(-1988, -3580);
        nextCycle(2383); checkResult(-1994, -3577);
        nextCycle(2384); checkResult(-1999, -3574);
        nextCycle(2385); checkResult(-2005, -3571);
        nextCycle(2386); checkResult(-2010, -3568);
        nextCycle(2387); checkResult(-2016, -3565);
        nextCycle(2388); checkResult(-2021, -3561);
        nextCycle(2389); checkResult(-2027, -3558);
        nextCycle(2390); checkResult(-2032, -3555);
        nextCycle(2391); checkResult(-2038, -3552);
        nextCycle(2392); checkResult(-2043, -3549);
        nextCycle(2393); checkResult(-2048, -3546);
        nextCycle(2394); checkResult(-2054, -3543);
        nextCycle(2395); checkResult(-2059, -3540);
        nextCycle(2396); checkResult(-2065, -3536);
        nextCycle(2397); checkResult(-2070, -3533);
        nextCycle(2398); checkResult(-2076, -3530);
        nextCycle(2399); checkResult(-2081, -3527);
        nextCycle(2400); checkResult(-2086, -3524);
        nextCycle(2401); checkResult(-2092, -3520);
        nextCycle(2402); checkResult(-2097, -3517);
        nextCycle(2403); checkResult(-2103, -3514);
        nextCycle(2404); checkResult(-2108, -3511);
        nextCycle(2405); checkResult(-2113, -3508);
        nextCycle(2406); checkResult(-2119, -3504);
        nextCycle(2407); checkResult(-2124, -3501);
        nextCycle(2408); checkResult(-2129, -3498);
        nextCycle(2409); checkResult(-2135, -3495);
        nextCycle(2410); checkResult(-2140, -3491);
        nextCycle(2411); checkResult(-2146, -3488);
        nextCycle(2412); checkResult(-2151, -3485);
        nextCycle(2413); checkResult(-2156, -3481);
        nextCycle(2414); checkResult(-2162, -3478);
        nextCycle(2415); checkResult(-2167, -3475);
        nextCycle(2416); checkResult(-2172, -3471);
        nextCycle(2417); checkResult(-2178, -3468);
        nextCycle(2418); checkResult(-2183, -3465);
        nextCycle(2419); checkResult(-2188, -3461);
        nextCycle(2420); checkResult(-2193, -3458);
        nextCycle(2421); checkResult(-2199, -3455);
        nextCycle(2422); checkResult(-2204, -3451);
        nextCycle(2423); checkResult(-2209, -3448);
        nextCycle(2424); checkResult(-2215, -3444);
        nextCycle(2425); checkResult(-2220, -3441);
        nextCycle(2426); checkResult(-2225, -3438);
        nextCycle(2427); checkResult(-2230, -3434);
        nextCycle(2428); checkResult(-2236, -3431);
        nextCycle(2429); checkResult(-2241, -3427);
        nextCycle(2430); checkResult(-2246, -3424);
        nextCycle(2431); checkResult(-2252, -3420);
        nextCycle(2432); checkResult(-2257, -3417);
        nextCycle(2433); checkResult(-2262, -3414);
        nextCycle(2434); checkResult(-2267, -3410);
        nextCycle(2435); checkResult(-2272, -3407);
        nextCycle(2436); checkResult(-2278, -3403);
        nextCycle(2437); checkResult(-2283, -3400);
        nextCycle(2438); checkResult(-2288, -3396);
        nextCycle(2439); checkResult(-2293, -3393);
        nextCycle(2440); checkResult(-2299, -3389);
        nextCycle(2441); checkResult(-2304, -3386);
        nextCycle(2442); checkResult(-2309, -3382);
        nextCycle(2443); checkResult(-2314, -3378);
        nextCycle(2444); checkResult(-2319, -3375);
        nextCycle(2445); checkResult(-2324, -3371);
        nextCycle(2446); checkResult(-2330, -3368);
        nextCycle(2447); checkResult(-2335, -3364);
        nextCycle(2448); checkResult(-2340, -3361);
        nextCycle(2449); checkResult(-2345, -3357);
        nextCycle(2450); checkResult(-2350, -3353);
        nextCycle(2451); checkResult(-2355, -3350);
        nextCycle(2452); checkResult(-2361, -3346);
        nextCycle(2453); checkResult(-2366, -3343);
        nextCycle(2454); checkResult(-2371, -3339);
        nextCycle(2455); checkResult(-2376, -3335);
        nextCycle(2456); checkResult(-2381, -3332);
        nextCycle(2457); checkResult(-2386, -3328);
        nextCycle(2458); checkResult(-2391, -3324);
        nextCycle(2459); checkResult(-2396, -3321);
        nextCycle(2460); checkResult(-2401, -3317);
        nextCycle(2461); checkResult(-2406, -3313);
        nextCycle(2462); checkResult(-2412, -3310);
        nextCycle(2463); checkResult(-2417, -3306);
        nextCycle(2464); checkResult(-2422, -3302);
        nextCycle(2465); checkResult(-2427, -3298);
        nextCycle(2466); checkResult(-2432, -3295);
        nextCycle(2467); checkResult(-2437, -3291);
        nextCycle(2468); checkResult(-2442, -3287);
        nextCycle(2469); checkResult(-2447, -3284);
        nextCycle(2470); checkResult(-2452, -3280);
        nextCycle(2471); checkResult(-2457, -3276);
        nextCycle(2472); checkResult(-2462, -3272);
        nextCycle(2473); checkResult(-2467, -3268);
        nextCycle(2474); checkResult(-2472, -3265);
        nextCycle(2475); checkResult(-2477, -3261);
        nextCycle(2476); checkResult(-2482, -3257);
        nextCycle(2477); checkResult(-2487, -3253);
        nextCycle(2478); checkResult(-2492, -3249);
        nextCycle(2479); checkResult(-2497, -3246);
        nextCycle(2480); checkResult(-2502, -3242);
        nextCycle(2481); checkResult(-2507, -3238);
        nextCycle(2482); checkResult(-2512, -3234);
        nextCycle(2483); checkResult(-2517, -3230);
        nextCycle(2484); checkResult(-2522, -3226);
        nextCycle(2485); checkResult(-2527, -3222);
        nextCycle(2486); checkResult(-2532, -3219);
        nextCycle(2487); checkResult(-2537, -3215);
        nextCycle(2488); checkResult(-2542, -3211);
        nextCycle(2489); checkResult(-2547, -3207);
        nextCycle(2490); checkResult(-2551, -3203);
        nextCycle(2491); checkResult(-2556, -3199);
        nextCycle(2492); checkResult(-2561, -3195);
        nextCycle(2493); checkResult(-2566, -3191);
        nextCycle(2494); checkResult(-2571, -3187);
        nextCycle(2495); checkResult(-2576, -3183);
        nextCycle(2496); checkResult(-2581, -3179);
        nextCycle(2497); checkResult(-2586, -3175);
        nextCycle(2498); checkResult(-2591, -3171);
        nextCycle(2499); checkResult(-2595, -3167);
        nextCycle(2500); checkResult(-2600, -3163);
        nextCycle(2501); checkResult(-2605, -3159);
        nextCycle(2502); checkResult(-2610, -3155);
        nextCycle(2503); checkResult(-2615, -3151);
        nextCycle(2504); checkResult(-2620, -3147);
        nextCycle(2505); checkResult(-2624, -3143);
        nextCycle(2506); checkResult(-2629, -3139);
        nextCycle(2507); checkResult(-2634, -3135);
        nextCycle(2508); checkResult(-2639, -3131);
        nextCycle(2509); checkResult(-2644, -3127);
        nextCycle(2510); checkResult(-2648, -3123);
        nextCycle(2511); checkResult(-2653, -3119);
        nextCycle(2512); checkResult(-2658, -3115);
        nextCycle(2513); checkResult(-2663, -3111);
        nextCycle(2514); checkResult(-2668, -3107);
        nextCycle(2515); checkResult(-2672, -3103);
        nextCycle(2516); checkResult(-2677, -3099);
        nextCycle(2517); checkResult(-2682, -3095);
        nextCycle(2518); checkResult(-2687, -3090);
        nextCycle(2519); checkResult(-2691, -3086);
        nextCycle(2520); checkResult(-2696, -3082);
        nextCycle(2521); checkResult(-2701, -3078);
        nextCycle(2522); checkResult(-2706, -3074);
        nextCycle(2523); checkResult(-2710, -3070);
        nextCycle(2524); checkResult(-2715, -3066);
        nextCycle(2525); checkResult(-2720, -3061);
        nextCycle(2526); checkResult(-2724, -3057);
        nextCycle(2527); checkResult(-2729, -3053);
        nextCycle(2528); checkResult(-2734, -3049);
        nextCycle(2529); checkResult(-2738, -3045);
        nextCycle(2530); checkResult(-2743, -3041);
        nextCycle(2531); checkResult(-2748, -3036);
        nextCycle(2532); checkResult(-2752, -3032);
        nextCycle(2533); checkResult(-2757, -3028);
        nextCycle(2534); checkResult(-2762, -3024);
        nextCycle(2535); checkResult(-2766, -3019);
        nextCycle(2536); checkResult(-2771, -3015);
        nextCycle(2537); checkResult(-2776, -3011);
        nextCycle(2538); checkResult(-2780, -3007);
        nextCycle(2539); checkResult(-2785, -3002);
        nextCycle(2540); checkResult(-2789, -2998);
        nextCycle(2541); checkResult(-2794, -2994);
        nextCycle(2542); checkResult(-2799, -2990);
        nextCycle(2543); checkResult(-2803, -2985);
        nextCycle(2544); checkResult(-2808, -2981);
        nextCycle(2545); checkResult(-2812, -2977);
        nextCycle(2546); checkResult(-2817, -2972);
        nextCycle(2547); checkResult(-2821, -2968);
        nextCycle(2548); checkResult(-2826, -2964);
        nextCycle(2549); checkResult(-2830, -2959);
        nextCycle(2550); checkResult(-2835, -2955);
        nextCycle(2551); checkResult(-2840, -2951);
        nextCycle(2552); checkResult(-2844, -2946);
        nextCycle(2553); checkResult(-2849, -2942);
        nextCycle(2554); checkResult(-2853, -2937);
        nextCycle(2555); checkResult(-2858, -2933);
        nextCycle(2556); checkResult(-2862, -2929);
        nextCycle(2557); checkResult(-2867, -2924);
        nextCycle(2558); checkResult(-2871, -2920);
        nextCycle(2559); checkResult(-2876, -2916);
        nextCycle(2560); checkResult(-2880, -2911);
        nextCycle(2561); checkResult(-2884, -2907);
        nextCycle(2562); checkResult(-2889, -2902);
        nextCycle(2563); checkResult(-2893, -2898);
        nextCycle(2564); checkResult(-2898, -2893);
        nextCycle(2565); checkResult(-2902, -2889);
        nextCycle(2566); checkResult(-2907, -2884);
        nextCycle(2567); checkResult(-2911, -2880);
        nextCycle(2568); checkResult(-2916, -2876);
        nextCycle(2569); checkResult(-2920, -2871);
        nextCycle(2570); checkResult(-2924, -2867);
        nextCycle(2571); checkResult(-2929, -2862);
        nextCycle(2572); checkResult(-2933, -2858);
        nextCycle(2573); checkResult(-2937, -2853);
        nextCycle(2574); checkResult(-2942, -2849);
        nextCycle(2575); checkResult(-2946, -2844);
        nextCycle(2576); checkResult(-2951, -2840);
        nextCycle(2577); checkResult(-2955, -2835);
        nextCycle(2578); checkResult(-2959, -2830);
        nextCycle(2579); checkResult(-2964, -2826);
        nextCycle(2580); checkResult(-2968, -2821);
        nextCycle(2581); checkResult(-2972, -2817);
        nextCycle(2582); checkResult(-2977, -2812);
        nextCycle(2583); checkResult(-2981, -2808);
        nextCycle(2584); checkResult(-2985, -2803);
        nextCycle(2585); checkResult(-2990, -2799);
        nextCycle(2586); checkResult(-2994, -2794);
        nextCycle(2587); checkResult(-2998, -2789);
        nextCycle(2588); checkResult(-3002, -2785);
        nextCycle(2589); checkResult(-3007, -2780);
        nextCycle(2590); checkResult(-3011, -2776);
        nextCycle(2591); checkResult(-3015, -2771);
        nextCycle(2592); checkResult(-3019, -2766);
        nextCycle(2593); checkResult(-3024, -2762);
        nextCycle(2594); checkResult(-3028, -2757);
        nextCycle(2595); checkResult(-3032, -2752);
        nextCycle(2596); checkResult(-3036, -2748);
        nextCycle(2597); checkResult(-3041, -2743);
        nextCycle(2598); checkResult(-3045, -2738);
        nextCycle(2599); checkResult(-3049, -2734);
        nextCycle(2600); checkResult(-3053, -2729);
        nextCycle(2601); checkResult(-3057, -2724);
        nextCycle(2602); checkResult(-3061, -2720);
        nextCycle(2603); checkResult(-3066, -2715);
        nextCycle(2604); checkResult(-3070, -2710);
        nextCycle(2605); checkResult(-3074, -2706);
        nextCycle(2606); checkResult(-3078, -2701);
        nextCycle(2607); checkResult(-3082, -2696);
        nextCycle(2608); checkResult(-3086, -2691);
        nextCycle(2609); checkResult(-3090, -2687);
        nextCycle(2610); checkResult(-3095, -2682);
        nextCycle(2611); checkResult(-3099, -2677);
        nextCycle(2612); checkResult(-3103, -2672);
        nextCycle(2613); checkResult(-3107, -2668);
        nextCycle(2614); checkResult(-3111, -2663);
        nextCycle(2615); checkResult(-3115, -2658);
        nextCycle(2616); checkResult(-3119, -2653);
        nextCycle(2617); checkResult(-3123, -2648);
        nextCycle(2618); checkResult(-3127, -2644);
        nextCycle(2619); checkResult(-3131, -2639);
        nextCycle(2620); checkResult(-3135, -2634);
        nextCycle(2621); checkResult(-3139, -2629);
        nextCycle(2622); checkResult(-3143, -2624);
        nextCycle(2623); checkResult(-3147, -2620);
        nextCycle(2624); checkResult(-3151, -2615);
        nextCycle(2625); checkResult(-3155, -2610);
        nextCycle(2626); checkResult(-3159, -2605);
        nextCycle(2627); checkResult(-3163, -2600);
        nextCycle(2628); checkResult(-3167, -2595);
        nextCycle(2629); checkResult(-3171, -2591);
        nextCycle(2630); checkResult(-3175, -2586);
        nextCycle(2631); checkResult(-3179, -2581);
        nextCycle(2632); checkResult(-3183, -2576);
        nextCycle(2633); checkResult(-3187, -2571);
        nextCycle(2634); checkResult(-3191, -2566);
        nextCycle(2635); checkResult(-3195, -2561);
        nextCycle(2636); checkResult(-3199, -2556);
        nextCycle(2637); checkResult(-3203, -2551);
        nextCycle(2638); checkResult(-3207, -2547);
        nextCycle(2639); checkResult(-3211, -2542);
        nextCycle(2640); checkResult(-3215, -2537);
        nextCycle(2641); checkResult(-3219, -2532);
        nextCycle(2642); checkResult(-3222, -2527);
        nextCycle(2643); checkResult(-3226, -2522);
        nextCycle(2644); checkResult(-3230, -2517);
        nextCycle(2645); checkResult(-3234, -2512);
        nextCycle(2646); checkResult(-3238, -2507);
        nextCycle(2647); checkResult(-3242, -2502);
        nextCycle(2648); checkResult(-3246, -2497);
        nextCycle(2649); checkResult(-3249, -2492);
        nextCycle(2650); checkResult(-3253, -2487);
        nextCycle(2651); checkResult(-3257, -2482);
        nextCycle(2652); checkResult(-3261, -2477);
        nextCycle(2653); checkResult(-3265, -2472);
        nextCycle(2654); checkResult(-3268, -2467);
        nextCycle(2655); checkResult(-3272, -2462);
        nextCycle(2656); checkResult(-3276, -2457);
        nextCycle(2657); checkResult(-3280, -2452);
        nextCycle(2658); checkResult(-3284, -2447);
        nextCycle(2659); checkResult(-3287, -2442);
        nextCycle(2660); checkResult(-3291, -2437);
        nextCycle(2661); checkResult(-3295, -2432);
        nextCycle(2662); checkResult(-3298, -2427);
        nextCycle(2663); checkResult(-3302, -2422);
        nextCycle(2664); checkResult(-3306, -2417);
        nextCycle(2665); checkResult(-3310, -2412);
        nextCycle(2666); checkResult(-3313, -2406);
        nextCycle(2667); checkResult(-3317, -2401);
        nextCycle(2668); checkResult(-3321, -2396);
        nextCycle(2669); checkResult(-3324, -2391);
        nextCycle(2670); checkResult(-3328, -2386);
        nextCycle(2671); checkResult(-3332, -2381);
        nextCycle(2672); checkResult(-3335, -2376);
        nextCycle(2673); checkResult(-3339, -2371);
        nextCycle(2674); checkResult(-3343, -2366);
        nextCycle(2675); checkResult(-3346, -2361);
        nextCycle(2676); checkResult(-3350, -2355);
        nextCycle(2677); checkResult(-3353, -2350);
        nextCycle(2678); checkResult(-3357, -2345);
        nextCycle(2679); checkResult(-3361, -2340);
        nextCycle(2680); checkResult(-3364, -2335);
        nextCycle(2681); checkResult(-3368, -2330);
        nextCycle(2682); checkResult(-3371, -2324);
        nextCycle(2683); checkResult(-3375, -2319);
        nextCycle(2684); checkResult(-3378, -2314);
        nextCycle(2685); checkResult(-3382, -2309);
        nextCycle(2686); checkResult(-3386, -2304);
        nextCycle(2687); checkResult(-3389, -2299);
        nextCycle(2688); checkResult(-3393, -2293);
        nextCycle(2689); checkResult(-3396, -2288);
        nextCycle(2690); checkResult(-3400, -2283);
        nextCycle(2691); checkResult(-3403, -2278);
        nextCycle(2692); checkResult(-3407, -2272);
        nextCycle(2693); checkResult(-3410, -2267);
        nextCycle(2694); checkResult(-3414, -2262);
        nextCycle(2695); checkResult(-3417, -2257);
        nextCycle(2696); checkResult(-3420, -2252);
        nextCycle(2697); checkResult(-3424, -2246);
        nextCycle(2698); checkResult(-3427, -2241);
        nextCycle(2699); checkResult(-3431, -2236);
        nextCycle(2700); checkResult(-3434, -2230);
        nextCycle(2701); checkResult(-3438, -2225);
        nextCycle(2702); checkResult(-3441, -2220);
        nextCycle(2703); checkResult(-3444, -2215);
        nextCycle(2704); checkResult(-3448, -2209);
        nextCycle(2705); checkResult(-3451, -2204);
        nextCycle(2706); checkResult(-3455, -2199);
        nextCycle(2707); checkResult(-3458, -2193);
        nextCycle(2708); checkResult(-3461, -2188);
        nextCycle(2709); checkResult(-3465, -2183);
        nextCycle(2710); checkResult(-3468, -2178);
        nextCycle(2711); checkResult(-3471, -2172);
        nextCycle(2712); checkResult(-3475, -2167);
        nextCycle(2713); checkResult(-3478, -2162);
        nextCycle(2714); checkResult(-3481, -2156);
        nextCycle(2715); checkResult(-3485, -2151);
        nextCycle(2716); checkResult(-3488, -2146);
        nextCycle(2717); checkResult(-3491, -2140);
        nextCycle(2718); checkResult(-3495, -2135);
        nextCycle(2719); checkResult(-3498, -2129);
        nextCycle(2720); checkResult(-3501, -2124);
        nextCycle(2721); checkResult(-3504, -2119);
        nextCycle(2722); checkResult(-3508, -2113);
        nextCycle(2723); checkResult(-3511, -2108);
        nextCycle(2724); checkResult(-3514, -2103);
        nextCycle(2725); checkResult(-3517, -2097);
        nextCycle(2726); checkResult(-3520, -2092);
        nextCycle(2727); checkResult(-3524, -2086);
        nextCycle(2728); checkResult(-3527, -2081);
        nextCycle(2729); checkResult(-3530, -2076);
        nextCycle(2730); checkResult(-3533, -2070);
        nextCycle(2731); checkResult(-3536, -2065);
        nextCycle(2732); checkResult(-3540, -2059);
        nextCycle(2733); checkResult(-3543, -2054);
        nextCycle(2734); checkResult(-3546, -2048);
        nextCycle(2735); checkResult(-3549, -2043);
        nextCycle(2736); checkResult(-3552, -2038);
        nextCycle(2737); checkResult(-3555, -2032);
        nextCycle(2738); checkResult(-3558, -2027);
        nextCycle(2739); checkResult(-3561, -2021);
        nextCycle(2740); checkResult(-3565, -2016);
        nextCycle(2741); checkResult(-3568, -2010);
        nextCycle(2742); checkResult(-3571, -2005);
        nextCycle(2743); checkResult(-3574, -1999);
        nextCycle(2744); checkResult(-3577, -1994);
        nextCycle(2745); checkResult(-3580, -1988);
        nextCycle(2746); checkResult(-3583, -1983);
        nextCycle(2747); checkResult(-3586, -1977);
        nextCycle(2748); checkResult(-3589, -1972);
        nextCycle(2749); checkResult(-3592, -1966);
        nextCycle(2750); checkResult(-3595, -1961);
        nextCycle(2751); checkResult(-3598, -1955);
        nextCycle(2752); checkResult(-3601, -1950);
        nextCycle(2753); checkResult(-3604, -1944);
        nextCycle(2754); checkResult(-3607, -1939);
        nextCycle(2755); checkResult(-3610, -1933);
        nextCycle(2756); checkResult(-3613, -1928);
        nextCycle(2757); checkResult(-3616, -1922);
        nextCycle(2758); checkResult(-3619, -1917);
        nextCycle(2759); checkResult(-3622, -1911);
        nextCycle(2760); checkResult(-3625, -1905);
        nextCycle(2761); checkResult(-3628, -1900);
        nextCycle(2762); checkResult(-3631, -1894);
        nextCycle(2763); checkResult(-3633, -1889);
        nextCycle(2764); checkResult(-3636, -1883);
        nextCycle(2765); checkResult(-3639, -1878);
        nextCycle(2766); checkResult(-3642, -1872);
        nextCycle(2767); checkResult(-3645, -1866);
        nextCycle(2768); checkResult(-3648, -1861);
        nextCycle(2769); checkResult(-3651, -1855);
        nextCycle(2770); checkResult(-3654, -1850);
        nextCycle(2771); checkResult(-3656, -1844);
        nextCycle(2772); checkResult(-3659, -1838);
        nextCycle(2773); checkResult(-3662, -1833);
        nextCycle(2774); checkResult(-3665, -1827);
        nextCycle(2775); checkResult(-3668, -1821);
        nextCycle(2776); checkResult(-3670, -1816);
        nextCycle(2777); checkResult(-3673, -1810);
        nextCycle(2778); checkResult(-3676, -1805);
        nextCycle(2779); checkResult(-3679, -1799);
        nextCycle(2780); checkResult(-3681, -1793);
        nextCycle(2781); checkResult(-3684, -1788);
        nextCycle(2782); checkResult(-3687, -1782);
        nextCycle(2783); checkResult(-3690, -1776);
        nextCycle(2784); checkResult(-3692, -1771);
        nextCycle(2785); checkResult(-3695, -1765);
        nextCycle(2786); checkResult(-3698, -1759);
        nextCycle(2787); checkResult(-3700, -1754);
        nextCycle(2788); checkResult(-3703, -1748);
        nextCycle(2789); checkResult(-3706, -1742);
        nextCycle(2790); checkResult(-3709, -1737);
        nextCycle(2791); checkResult(-3711, -1731);
        nextCycle(2792); checkResult(-3714, -1725);
        nextCycle(2793); checkResult(-3716, -1720);
        nextCycle(2794); checkResult(-3719, -1714);
        nextCycle(2795); checkResult(-3722, -1708);
        nextCycle(2796); checkResult(-3724, -1702);
        nextCycle(2797); checkResult(-3727, -1697);
        nextCycle(2798); checkResult(-3730, -1691);
        nextCycle(2799); checkResult(-3732, -1685);
        nextCycle(2800); checkResult(-3735, -1680);
        nextCycle(2801); checkResult(-3737, -1674);
        nextCycle(2802); checkResult(-3740, -1668);
        nextCycle(2803); checkResult(-3742, -1662);
        nextCycle(2804); checkResult(-3745, -1657);
        nextCycle(2805); checkResult(-3747, -1651);
        nextCycle(2806); checkResult(-3750, -1645);
        nextCycle(2807); checkResult(-3753, -1639);
        nextCycle(2808); checkResult(-3755, -1634);
        nextCycle(2809); checkResult(-3758, -1628);
        nextCycle(2810); checkResult(-3760, -1622);
        nextCycle(2811); checkResult(-3763, -1616);
        nextCycle(2812); checkResult(-3765, -1611);
        nextCycle(2813); checkResult(-3767, -1605);
        nextCycle(2814); checkResult(-3770, -1599);
        nextCycle(2815); checkResult(-3772, -1593);
        nextCycle(2816); checkResult(-3775, -1587);
        nextCycle(2817); checkResult(-3777, -1582);
        nextCycle(2818); checkResult(-3780, -1576);
        nextCycle(2819); checkResult(-3782, -1570);
        nextCycle(2820); checkResult(-3784, -1564);
        nextCycle(2821); checkResult(-3787, -1558);
        nextCycle(2822); checkResult(-3789, -1553);
        nextCycle(2823); checkResult(-3792, -1547);
        nextCycle(2824); checkResult(-3794, -1541);
        nextCycle(2825); checkResult(-3796, -1535);
        nextCycle(2826); checkResult(-3799, -1529);
        nextCycle(2827); checkResult(-3801, -1523);
        nextCycle(2828); checkResult(-3803, -1518);
        nextCycle(2829); checkResult(-3806, -1512);
        nextCycle(2830); checkResult(-3808, -1506);
        nextCycle(2831); checkResult(-3810, -1500);
        nextCycle(2832); checkResult(-3813, -1494);
        nextCycle(2833); checkResult(-3815, -1488);
        nextCycle(2834); checkResult(-3817, -1483);
        nextCycle(2835); checkResult(-3819, -1477);
        nextCycle(2836); checkResult(-3822, -1471);
        nextCycle(2837); checkResult(-3824, -1465);
        nextCycle(2838); checkResult(-3826, -1459);
        nextCycle(2839); checkResult(-3828, -1453);
        nextCycle(2840); checkResult(-3831, -1447);
        nextCycle(2841); checkResult(-3833, -1441);
        nextCycle(2842); checkResult(-3835, -1436);
        nextCycle(2843); checkResult(-3837, -1430);
        nextCycle(2844); checkResult(-3839, -1424);
        nextCycle(2845); checkResult(-3842, -1418);
        nextCycle(2846); checkResult(-3844, -1412);
        nextCycle(2847); checkResult(-3846, -1406);
        nextCycle(2848); checkResult(-3848, -1400);
        nextCycle(2849); checkResult(-3850, -1394);
        nextCycle(2850); checkResult(-3852, -1388);
        nextCycle(2851); checkResult(-3855, -1383);
        nextCycle(2852); checkResult(-3857, -1377);
        nextCycle(2853); checkResult(-3859, -1371);
        nextCycle(2854); checkResult(-3861, -1365);
        nextCycle(2855); checkResult(-3863, -1359);
        nextCycle(2856); checkResult(-3865, -1353);
        nextCycle(2857); checkResult(-3867, -1347);
        nextCycle(2858); checkResult(-3869, -1341);
        nextCycle(2859); checkResult(-3871, -1335);
        nextCycle(2860); checkResult(-3873, -1329);
        nextCycle(2861); checkResult(-3875, -1323);
        nextCycle(2862); checkResult(-3877, -1317);
        nextCycle(2863); checkResult(-3879, -1311);
        nextCycle(2864); checkResult(-3881, -1305);
        nextCycle(2865); checkResult(-3883, -1299);
        nextCycle(2866); checkResult(-3885, -1293);
        nextCycle(2867); checkResult(-3887, -1288);
        nextCycle(2868); checkResult(-3889, -1282);
        nextCycle(2869); checkResult(-3891, -1276);
        nextCycle(2870); checkResult(-3893, -1270);
        nextCycle(2871); checkResult(-3895, -1264);
        nextCycle(2872); checkResult(-3897, -1258);
        nextCycle(2873); checkResult(-3899, -1252);
        nextCycle(2874); checkResult(-3901, -1246);
        nextCycle(2875); checkResult(-3903, -1240);
        nextCycle(2876); checkResult(-3905, -1234);
        nextCycle(2877); checkResult(-3907, -1228);
        nextCycle(2878); checkResult(-3909, -1222);
        nextCycle(2879); checkResult(-3910, -1216);
        nextCycle(2880); checkResult(-3912, -1210);
        nextCycle(2881); checkResult(-3914, -1204);
        nextCycle(2882); checkResult(-3916, -1198);
        nextCycle(2883); checkResult(-3918, -1192);
        nextCycle(2884); checkResult(-3920, -1186);
        nextCycle(2885); checkResult(-3921, -1180);
        nextCycle(2886); checkResult(-3923, -1174);
        nextCycle(2887); checkResult(-3925, -1168);
        nextCycle(2888); checkResult(-3927, -1162);
        nextCycle(2889); checkResult(-3929, -1156);
        nextCycle(2890); checkResult(-3930, -1150);
        nextCycle(2891); checkResult(-3932, -1144);
        nextCycle(2892); checkResult(-3934, -1138);
        nextCycle(2893); checkResult(-3936, -1131);
        nextCycle(2894); checkResult(-3937, -1125);
        nextCycle(2895); checkResult(-3939, -1119);
        nextCycle(2896); checkResult(-3941, -1113);
        nextCycle(2897); checkResult(-3942, -1107);
        nextCycle(2898); checkResult(-3944, -1101);
        nextCycle(2899); checkResult(-3946, -1095);
        nextCycle(2900); checkResult(-3947, -1089);
        nextCycle(2901); checkResult(-3949, -1083);
        nextCycle(2902); checkResult(-3951, -1077);
        nextCycle(2903); checkResult(-3952, -1071);
        nextCycle(2904); checkResult(-3954, -1065);
        nextCycle(2905); checkResult(-3956, -1059);
        nextCycle(2906); checkResult(-3957, -1053);
        nextCycle(2907); checkResult(-3959, -1047);
        nextCycle(2908); checkResult(-3961, -1041);
        nextCycle(2909); checkResult(-3962, -1035);
        nextCycle(2910); checkResult(-3964, -1028);
        nextCycle(2911); checkResult(-3965, -1022);
        nextCycle(2912); checkResult(-3967, -1016);
        nextCycle(2913); checkResult(-3968, -1010);
        nextCycle(2914); checkResult(-3970, -1004);
        nextCycle(2915); checkResult(-3972, -998);
        nextCycle(2916); checkResult(-3973, -992);
        nextCycle(2917); checkResult(-3975, -986);
        nextCycle(2918); checkResult(-3976, -980);
        nextCycle(2919); checkResult(-3978, -974);
        nextCycle(2920); checkResult(-3979, -968);
        nextCycle(2921); checkResult(-3981, -961);
        nextCycle(2922); checkResult(-3982, -955);
        nextCycle(2923); checkResult(-3983, -949);
        nextCycle(2924); checkResult(-3985, -943);
        nextCycle(2925); checkResult(-3986, -937);
        nextCycle(2926); checkResult(-3988, -931);
        nextCycle(2927); checkResult(-3989, -925);
        nextCycle(2928); checkResult(-3991, -919);
        nextCycle(2929); checkResult(-3992, -913);
        nextCycle(2930); checkResult(-3993, -906);
        nextCycle(2931); checkResult(-3995, -900);
        nextCycle(2932); checkResult(-3996, -894);
        nextCycle(2933); checkResult(-3998, -888);
        nextCycle(2934); checkResult(-3999, -882);
        nextCycle(2935); checkResult(-4000, -876);
        nextCycle(2936); checkResult(-4002, -870);
        nextCycle(2937); checkResult(-4003, -863);
        nextCycle(2938); checkResult(-4004, -857);
        nextCycle(2939); checkResult(-4006, -851);
        nextCycle(2940); checkResult(-4007, -845);
        nextCycle(2941); checkResult(-4008, -839);
        nextCycle(2942); checkResult(-4009, -833);
        nextCycle(2943); checkResult(-4011, -827);
        nextCycle(2944); checkResult(-4012, -820);
        nextCycle(2945); checkResult(-4013, -814);
        nextCycle(2946); checkResult(-4014, -808);
        nextCycle(2947); checkResult(-4016, -802);
        nextCycle(2948); checkResult(-4017, -796);
        nextCycle(2949); checkResult(-4018, -790);
        nextCycle(2950); checkResult(-4019, -783);
        nextCycle(2951); checkResult(-4021, -777);
        nextCycle(2952); checkResult(-4022, -771);
        nextCycle(2953); checkResult(-4023, -765);
        nextCycle(2954); checkResult(-4024, -759);
        nextCycle(2955); checkResult(-4025, -753);
        nextCycle(2956); checkResult(-4026, -746);
        nextCycle(2957); checkResult(-4028, -740);
        nextCycle(2958); checkResult(-4029, -734);
        nextCycle(2959); checkResult(-4030, -728);
        nextCycle(2960); checkResult(-4031, -722);
        nextCycle(2961); checkResult(-4032, -716);
        nextCycle(2962); checkResult(-4033, -709);
        nextCycle(2963); checkResult(-4034, -703);
        nextCycle(2964); checkResult(-4035, -697);
        nextCycle(2965); checkResult(-4036, -691);
        nextCycle(2966); checkResult(-4037, -685);
        nextCycle(2967); checkResult(-4038, -678);
        nextCycle(2968); checkResult(-4039, -672);
        nextCycle(2969); checkResult(-4040, -666);
        nextCycle(2970); checkResult(-4041, -660);
        nextCycle(2971); checkResult(-4042, -654);
        nextCycle(2972); checkResult(-4043, -647);
        nextCycle(2973); checkResult(-4044, -641);
        nextCycle(2974); checkResult(-4045, -635);
        nextCycle(2975); checkResult(-4046, -629);
        nextCycle(2976); checkResult(-4047, -623);
        nextCycle(2977); checkResult(-4048, -616);
        nextCycle(2978); checkResult(-4049, -610);
        nextCycle(2979); checkResult(-4050, -604);
        nextCycle(2980); checkResult(-4051, -598);
        nextCycle(2981); checkResult(-4052, -592);
        nextCycle(2982); checkResult(-4053, -585);
        nextCycle(2983); checkResult(-4054, -579);
        nextCycle(2984); checkResult(-4055, -573);
        nextCycle(2985); checkResult(-4056, -567);
        nextCycle(2986); checkResult(-4056, -560);
        nextCycle(2987); checkResult(-4057, -554);
        nextCycle(2988); checkResult(-4058, -548);
        nextCycle(2989); checkResult(-4059, -542);
        nextCycle(2990); checkResult(-4060, -536);
        nextCycle(2991); checkResult(-4061, -529);
        nextCycle(2992); checkResult(-4061, -523);
        nextCycle(2993); checkResult(-4062, -517);
        nextCycle(2994); checkResult(-4063, -511);
        nextCycle(2995); checkResult(-4064, -504);
        nextCycle(2996); checkResult(-4065, -498);
        nextCycle(2997); checkResult(-4065, -492);
        nextCycle(2998); checkResult(-4066, -486);
        nextCycle(2999); checkResult(-4067, -479);
        nextCycle(3000); checkResult(-4068, -473);
        nextCycle(3001); checkResult(-4068, -467);
        nextCycle(3002); checkResult(-4069, -461);
        nextCycle(3003); checkResult(-4070, -454);
        nextCycle(3004); checkResult(-4070, -448);
        nextCycle(3005); checkResult(-4071, -442);
        nextCycle(3006); checkResult(-4072, -436);
        nextCycle(3007); checkResult(-4072, -430);
        nextCycle(3008); checkResult(-4073, -423);
        nextCycle(3009); checkResult(-4074, -417);
        nextCycle(3010); checkResult(-4074, -411);
        nextCycle(3011); checkResult(-4075, -405);
        nextCycle(3012); checkResult(-4076, -398);
        nextCycle(3013); checkResult(-4076, -392);
        nextCycle(3014); checkResult(-4077, -386);
        nextCycle(3015); checkResult(-4077, -379);
        nextCycle(3016); checkResult(-4078, -373);
        nextCycle(3017); checkResult(-4079, -367);
        nextCycle(3018); checkResult(-4079, -361);
        nextCycle(3019); checkResult(-4080, -354);
        nextCycle(3020); checkResult(-4080, -348);
        nextCycle(3021); checkResult(-4081, -342);
        nextCycle(3022); checkResult(-4081, -336);
        nextCycle(3023); checkResult(-4082, -329);
        nextCycle(3024); checkResult(-4082, -323);
        nextCycle(3025); checkResult(-4083, -317);
        nextCycle(3026); checkResult(-4083, -311);
        nextCycle(3027); checkResult(-4084, -304);
        nextCycle(3028); checkResult(-4084, -298);
        nextCycle(3029); checkResult(-4085, -292);
        nextCycle(3030); checkResult(-4085, -286);
        nextCycle(3031); checkResult(-4085, -279);
        nextCycle(3032); checkResult(-4086, -273);
        nextCycle(3033); checkResult(-4086, -267);
        nextCycle(3034); checkResult(-4087, -261);
        nextCycle(3035); checkResult(-4087, -254);
        nextCycle(3036); checkResult(-4087, -248);
        nextCycle(3037); checkResult(-4088, -242);
        nextCycle(3038); checkResult(-4088, -235);
        nextCycle(3039); checkResult(-4089, -229);
        nextCycle(3040); checkResult(-4089, -223);
        nextCycle(3041); checkResult(-4089, -217);
        nextCycle(3042); checkResult(-4090, -210);
        nextCycle(3043); checkResult(-4090, -204);
        nextCycle(3044); checkResult(-4090, -198);
        nextCycle(3045); checkResult(-4091, -192);
        nextCycle(3046); checkResult(-4091, -185);
        nextCycle(3047); checkResult(-4091, -179);
        nextCycle(3048); checkResult(-4091, -173);
        nextCycle(3049); checkResult(-4092, -166);
        nextCycle(3050); checkResult(-4092, -160);
        nextCycle(3051); checkResult(-4092, -154);
        nextCycle(3052); checkResult(-4092, -148);
        nextCycle(3053); checkResult(-4093, -141);
        nextCycle(3054); checkResult(-4093, -135);
        nextCycle(3055); checkResult(-4093, -129);
        nextCycle(3056); checkResult(-4093, -122);
        nextCycle(3057); checkResult(-4093, -116);
        nextCycle(3058); checkResult(-4094, -110);
        nextCycle(3059); checkResult(-4094, -104);
        nextCycle(3060); checkResult(-4094, -97);
        nextCycle(3061); checkResult(-4094, -91);
        nextCycle(3062); checkResult(-4094, -85);
        nextCycle(3063); checkResult(-4094, -79);
        nextCycle(3064); checkResult(-4094, -72);
        nextCycle(3065); checkResult(-4094, -66);
        nextCycle(3066); checkResult(-4095, -60);
        nextCycle(3067); checkResult(-4095, -53);
        nextCycle(3068); checkResult(-4095, -47);
        nextCycle(3069); checkResult(-4095, -41);
        nextCycle(3070); checkResult(-4095, -35);
        nextCycle(3071); checkResult(-4095, -28);
        nextCycle(3072); checkResult(-4095, -22);
        nextCycle(3073); checkResult(-4095, -16);
        nextCycle(3074); checkResult(-4095, -9);
        nextCycle(3075); checkResult(-4095, -3);
        nextCycle(3076); checkResult(-4095, 3);
        nextCycle(3077); checkResult(-4095, 9);
        nextCycle(3078); checkResult(-4095, 16);
        nextCycle(3079); checkResult(-4095, 22);
        nextCycle(3080); checkResult(-4095, 28);
        nextCycle(3081); checkResult(-4095, 35);
        nextCycle(3082); checkResult(-4095, 41);
        nextCycle(3083); checkResult(-4095, 47);
        nextCycle(3084); checkResult(-4095, 53);
        nextCycle(3085); checkResult(-4095, 60);
        nextCycle(3086); checkResult(-4094, 66);
        nextCycle(3087); checkResult(-4094, 72);
        nextCycle(3088); checkResult(-4094, 79);
        nextCycle(3089); checkResult(-4094, 85);
        nextCycle(3090); checkResult(-4094, 91);
        nextCycle(3091); checkResult(-4094, 97);
        nextCycle(3092); checkResult(-4094, 104);
        nextCycle(3093); checkResult(-4094, 110);
        nextCycle(3094); checkResult(-4093, 116);
        nextCycle(3095); checkResult(-4093, 122);
        nextCycle(3096); checkResult(-4093, 129);
        nextCycle(3097); checkResult(-4093, 135);
        nextCycle(3098); checkResult(-4093, 141);
        nextCycle(3099); checkResult(-4092, 148);
        nextCycle(3100); checkResult(-4092, 154);
        nextCycle(3101); checkResult(-4092, 160);
        nextCycle(3102); checkResult(-4092, 166);
        nextCycle(3103); checkResult(-4091, 173);
        nextCycle(3104); checkResult(-4091, 179);
        nextCycle(3105); checkResult(-4091, 185);
        nextCycle(3106); checkResult(-4091, 192);
        nextCycle(3107); checkResult(-4090, 198);
        nextCycle(3108); checkResult(-4090, 204);
        nextCycle(3109); checkResult(-4090, 210);
        nextCycle(3110); checkResult(-4089, 217);
        nextCycle(3111); checkResult(-4089, 223);
        nextCycle(3112); checkResult(-4089, 229);
        nextCycle(3113); checkResult(-4088, 235);
        nextCycle(3114); checkResult(-4088, 242);
        nextCycle(3115); checkResult(-4087, 248);
        nextCycle(3116); checkResult(-4087, 254);
        nextCycle(3117); checkResult(-4087, 261);
        nextCycle(3118); checkResult(-4086, 267);
        nextCycle(3119); checkResult(-4086, 273);
        nextCycle(3120); checkResult(-4085, 279);
        nextCycle(3121); checkResult(-4085, 286);
        nextCycle(3122); checkResult(-4085, 292);
        nextCycle(3123); checkResult(-4084, 298);
        nextCycle(3124); checkResult(-4084, 304);
        nextCycle(3125); checkResult(-4083, 311);
        nextCycle(3126); checkResult(-4083, 317);
        nextCycle(3127); checkResult(-4082, 323);
        nextCycle(3128); checkResult(-4082, 329);
        nextCycle(3129); checkResult(-4081, 336);
        nextCycle(3130); checkResult(-4081, 342);
        nextCycle(3131); checkResult(-4080, 348);
        nextCycle(3132); checkResult(-4080, 354);
        nextCycle(3133); checkResult(-4079, 361);
        nextCycle(3134); checkResult(-4079, 367);
        nextCycle(3135); checkResult(-4078, 373);
        nextCycle(3136); checkResult(-4077, 379);
        nextCycle(3137); checkResult(-4077, 386);
        nextCycle(3138); checkResult(-4076, 392);
        nextCycle(3139); checkResult(-4076, 398);
        nextCycle(3140); checkResult(-4075, 405);
        nextCycle(3141); checkResult(-4074, 411);
        nextCycle(3142); checkResult(-4074, 417);
        nextCycle(3143); checkResult(-4073, 423);
        nextCycle(3144); checkResult(-4072, 430);
        nextCycle(3145); checkResult(-4072, 436);
        nextCycle(3146); checkResult(-4071, 442);
        nextCycle(3147); checkResult(-4070, 448);
        nextCycle(3148); checkResult(-4070, 454);
        nextCycle(3149); checkResult(-4069, 461);
        nextCycle(3150); checkResult(-4068, 467);
        nextCycle(3151); checkResult(-4068, 473);
        nextCycle(3152); checkResult(-4067, 479);
        nextCycle(3153); checkResult(-4066, 486);
        nextCycle(3154); checkResult(-4065, 492);
        nextCycle(3155); checkResult(-4065, 498);
        nextCycle(3156); checkResult(-4064, 504);
        nextCycle(3157); checkResult(-4063, 511);
        nextCycle(3158); checkResult(-4062, 517);
        nextCycle(3159); checkResult(-4061, 523);
        nextCycle(3160); checkResult(-4061, 529);
        nextCycle(3161); checkResult(-4060, 536);
        nextCycle(3162); checkResult(-4059, 542);
        nextCycle(3163); checkResult(-4058, 548);
        nextCycle(3164); checkResult(-4057, 554);
        nextCycle(3165); checkResult(-4056, 560);
        nextCycle(3166); checkResult(-4056, 567);
        nextCycle(3167); checkResult(-4055, 573);
        nextCycle(3168); checkResult(-4054, 579);
        nextCycle(3169); checkResult(-4053, 585);
        nextCycle(3170); checkResult(-4052, 592);
        nextCycle(3171); checkResult(-4051, 598);
        nextCycle(3172); checkResult(-4050, 604);
        nextCycle(3173); checkResult(-4049, 610);
        nextCycle(3174); checkResult(-4048, 616);
        nextCycle(3175); checkResult(-4047, 623);
        nextCycle(3176); checkResult(-4046, 629);
        nextCycle(3177); checkResult(-4045, 635);
        nextCycle(3178); checkResult(-4044, 641);
        nextCycle(3179); checkResult(-4043, 647);
        nextCycle(3180); checkResult(-4042, 654);
        nextCycle(3181); checkResult(-4041, 660);
        nextCycle(3182); checkResult(-4040, 666);
        nextCycle(3183); checkResult(-4039, 672);
        nextCycle(3184); checkResult(-4038, 678);
        nextCycle(3185); checkResult(-4037, 685);
        nextCycle(3186); checkResult(-4036, 691);
        nextCycle(3187); checkResult(-4035, 697);
        nextCycle(3188); checkResult(-4034, 703);
        nextCycle(3189); checkResult(-4033, 709);
        nextCycle(3190); checkResult(-4032, 716);
        nextCycle(3191); checkResult(-4031, 722);
        nextCycle(3192); checkResult(-4030, 728);
        nextCycle(3193); checkResult(-4029, 734);
        nextCycle(3194); checkResult(-4028, 740);
        nextCycle(3195); checkResult(-4026, 746);
        nextCycle(3196); checkResult(-4025, 753);
        nextCycle(3197); checkResult(-4024, 759);
        nextCycle(3198); checkResult(-4023, 765);
        nextCycle(3199); checkResult(-4022, 771);
        nextCycle(3200); checkResult(-4021, 777);
        nextCycle(3201); checkResult(-4019, 783);
        nextCycle(3202); checkResult(-4018, 790);
        nextCycle(3203); checkResult(-4017, 796);
        nextCycle(3204); checkResult(-4016, 802);
        nextCycle(3205); checkResult(-4014, 808);
        nextCycle(3206); checkResult(-4013, 814);
        nextCycle(3207); checkResult(-4012, 820);
        nextCycle(3208); checkResult(-4011, 827);
        nextCycle(3209); checkResult(-4009, 833);
        nextCycle(3210); checkResult(-4008, 839);
        nextCycle(3211); checkResult(-4007, 845);
        nextCycle(3212); checkResult(-4006, 851);
        nextCycle(3213); checkResult(-4004, 857);
        nextCycle(3214); checkResult(-4003, 863);
        nextCycle(3215); checkResult(-4002, 870);
        nextCycle(3216); checkResult(-4000, 876);
        nextCycle(3217); checkResult(-3999, 882);
        nextCycle(3218); checkResult(-3998, 888);
        nextCycle(3219); checkResult(-3996, 894);
        nextCycle(3220); checkResult(-3995, 900);
        nextCycle(3221); checkResult(-3993, 906);
        nextCycle(3222); checkResult(-3992, 913);
        nextCycle(3223); checkResult(-3991, 919);
        nextCycle(3224); checkResult(-3989, 925);
        nextCycle(3225); checkResult(-3988, 931);
        nextCycle(3226); checkResult(-3986, 937);
        nextCycle(3227); checkResult(-3985, 943);
        nextCycle(3228); checkResult(-3983, 949);
        nextCycle(3229); checkResult(-3982, 955);
        nextCycle(3230); checkResult(-3981, 961);
        nextCycle(3231); checkResult(-3979, 968);
        nextCycle(3232); checkResult(-3978, 974);
        nextCycle(3233); checkResult(-3976, 980);
        nextCycle(3234); checkResult(-3975, 986);
        nextCycle(3235); checkResult(-3973, 992);
        nextCycle(3236); checkResult(-3972, 998);
        nextCycle(3237); checkResult(-3970, 1004);
        nextCycle(3238); checkResult(-3968, 1010);
        nextCycle(3239); checkResult(-3967, 1016);
        nextCycle(3240); checkResult(-3965, 1022);
        nextCycle(3241); checkResult(-3964, 1028);
        nextCycle(3242); checkResult(-3962, 1035);
        nextCycle(3243); checkResult(-3961, 1041);
        nextCycle(3244); checkResult(-3959, 1047);
        nextCycle(3245); checkResult(-3957, 1053);
        nextCycle(3246); checkResult(-3956, 1059);
        nextCycle(3247); checkResult(-3954, 1065);
        nextCycle(3248); checkResult(-3952, 1071);
        nextCycle(3249); checkResult(-3951, 1077);
        nextCycle(3250); checkResult(-3949, 1083);
        nextCycle(3251); checkResult(-3947, 1089);
        nextCycle(3252); checkResult(-3946, 1095);
        nextCycle(3253); checkResult(-3944, 1101);
        nextCycle(3254); checkResult(-3942, 1107);
        nextCycle(3255); checkResult(-3941, 1113);
        nextCycle(3256); checkResult(-3939, 1119);
        nextCycle(3257); checkResult(-3937, 1125);
        nextCycle(3258); checkResult(-3936, 1131);
        nextCycle(3259); checkResult(-3934, 1138);
        nextCycle(3260); checkResult(-3932, 1144);
        nextCycle(3261); checkResult(-3930, 1150);
        nextCycle(3262); checkResult(-3929, 1156);
        nextCycle(3263); checkResult(-3927, 1162);
        nextCycle(3264); checkResult(-3925, 1168);
        nextCycle(3265); checkResult(-3923, 1174);
        nextCycle(3266); checkResult(-3921, 1180);
        nextCycle(3267); checkResult(-3920, 1186);
        nextCycle(3268); checkResult(-3918, 1192);
        nextCycle(3269); checkResult(-3916, 1198);
        nextCycle(3270); checkResult(-3914, 1204);
        nextCycle(3271); checkResult(-3912, 1210);
        nextCycle(3272); checkResult(-3910, 1216);
        nextCycle(3273); checkResult(-3909, 1222);
        nextCycle(3274); checkResult(-3907, 1228);
        nextCycle(3275); checkResult(-3905, 1234);
        nextCycle(3276); checkResult(-3903, 1240);
        nextCycle(3277); checkResult(-3901, 1246);
        nextCycle(3278); checkResult(-3899, 1252);
        nextCycle(3279); checkResult(-3897, 1258);
        nextCycle(3280); checkResult(-3895, 1264);
        nextCycle(3281); checkResult(-3893, 1270);
        nextCycle(3282); checkResult(-3891, 1276);
        nextCycle(3283); checkResult(-3889, 1282);
        nextCycle(3284); checkResult(-3887, 1288);
        nextCycle(3285); checkResult(-3885, 1293);
        nextCycle(3286); checkResult(-3883, 1299);
        nextCycle(3287); checkResult(-3881, 1305);
        nextCycle(3288); checkResult(-3879, 1311);
        nextCycle(3289); checkResult(-3877, 1317);
        nextCycle(3290); checkResult(-3875, 1323);
        nextCycle(3291); checkResult(-3873, 1329);
        nextCycle(3292); checkResult(-3871, 1335);
        nextCycle(3293); checkResult(-3869, 1341);
        nextCycle(3294); checkResult(-3867, 1347);
        nextCycle(3295); checkResult(-3865, 1353);
        nextCycle(3296); checkResult(-3863, 1359);
        nextCycle(3297); checkResult(-3861, 1365);
        nextCycle(3298); checkResult(-3859, 1371);
        nextCycle(3299); checkResult(-3857, 1377);
        nextCycle(3300); checkResult(-3855, 1383);
        nextCycle(3301); checkResult(-3852, 1388);
        nextCycle(3302); checkResult(-3850, 1394);
        nextCycle(3303); checkResult(-3848, 1400);
        nextCycle(3304); checkResult(-3846, 1406);
        nextCycle(3305); checkResult(-3844, 1412);
        nextCycle(3306); checkResult(-3842, 1418);
        nextCycle(3307); checkResult(-3839, 1424);
        nextCycle(3308); checkResult(-3837, 1430);
        nextCycle(3309); checkResult(-3835, 1436);
        nextCycle(3310); checkResult(-3833, 1441);
        nextCycle(3311); checkResult(-3831, 1447);
        nextCycle(3312); checkResult(-3828, 1453);
        nextCycle(3313); checkResult(-3826, 1459);
        nextCycle(3314); checkResult(-3824, 1465);
        nextCycle(3315); checkResult(-3822, 1471);
        nextCycle(3316); checkResult(-3819, 1477);
        nextCycle(3317); checkResult(-3817, 1483);
        nextCycle(3318); checkResult(-3815, 1488);
        nextCycle(3319); checkResult(-3813, 1494);
        nextCycle(3320); checkResult(-3810, 1500);
        nextCycle(3321); checkResult(-3808, 1506);
        nextCycle(3322); checkResult(-3806, 1512);
        nextCycle(3323); checkResult(-3803, 1518);
        nextCycle(3324); checkResult(-3801, 1523);
        nextCycle(3325); checkResult(-3799, 1529);
        nextCycle(3326); checkResult(-3796, 1535);
        nextCycle(3327); checkResult(-3794, 1541);
        nextCycle(3328); checkResult(-3792, 1547);
        nextCycle(3329); checkResult(-3789, 1553);
        nextCycle(3330); checkResult(-3787, 1558);
        nextCycle(3331); checkResult(-3784, 1564);
        nextCycle(3332); checkResult(-3782, 1570);
        nextCycle(3333); checkResult(-3780, 1576);
        nextCycle(3334); checkResult(-3777, 1582);
        nextCycle(3335); checkResult(-3775, 1587);
        nextCycle(3336); checkResult(-3772, 1593);
        nextCycle(3337); checkResult(-3770, 1599);
        nextCycle(3338); checkResult(-3767, 1605);
        nextCycle(3339); checkResult(-3765, 1611);
        nextCycle(3340); checkResult(-3763, 1616);
        nextCycle(3341); checkResult(-3760, 1622);
        nextCycle(3342); checkResult(-3758, 1628);
        nextCycle(3343); checkResult(-3755, 1634);
        nextCycle(3344); checkResult(-3753, 1639);
        nextCycle(3345); checkResult(-3750, 1645);
        nextCycle(3346); checkResult(-3747, 1651);
        nextCycle(3347); checkResult(-3745, 1657);
        nextCycle(3348); checkResult(-3742, 1662);
        nextCycle(3349); checkResult(-3740, 1668);
        nextCycle(3350); checkResult(-3737, 1674);
        nextCycle(3351); checkResult(-3735, 1680);
        nextCycle(3352); checkResult(-3732, 1685);
        nextCycle(3353); checkResult(-3730, 1691);
        nextCycle(3354); checkResult(-3727, 1697);
        nextCycle(3355); checkResult(-3724, 1702);
        nextCycle(3356); checkResult(-3722, 1708);
        nextCycle(3357); checkResult(-3719, 1714);
        nextCycle(3358); checkResult(-3716, 1720);
        nextCycle(3359); checkResult(-3714, 1725);
        nextCycle(3360); checkResult(-3711, 1731);
        nextCycle(3361); checkResult(-3709, 1737);
        nextCycle(3362); checkResult(-3706, 1742);
        nextCycle(3363); checkResult(-3703, 1748);
        nextCycle(3364); checkResult(-3700, 1754);
        nextCycle(3365); checkResult(-3698, 1759);
        nextCycle(3366); checkResult(-3695, 1765);
        nextCycle(3367); checkResult(-3692, 1771);
        nextCycle(3368); checkResult(-3690, 1776);
        nextCycle(3369); checkResult(-3687, 1782);
        nextCycle(3370); checkResult(-3684, 1788);
        nextCycle(3371); checkResult(-3681, 1793);
        nextCycle(3372); checkResult(-3679, 1799);
        nextCycle(3373); checkResult(-3676, 1805);
        nextCycle(3374); checkResult(-3673, 1810);
        nextCycle(3375); checkResult(-3670, 1816);
        nextCycle(3376); checkResult(-3668, 1821);
        nextCycle(3377); checkResult(-3665, 1827);
        nextCycle(3378); checkResult(-3662, 1833);
        nextCycle(3379); checkResult(-3659, 1838);
        nextCycle(3380); checkResult(-3656, 1844);
        nextCycle(3381); checkResult(-3654, 1850);
        nextCycle(3382); checkResult(-3651, 1855);
        nextCycle(3383); checkResult(-3648, 1861);
        nextCycle(3384); checkResult(-3645, 1866);
        nextCycle(3385); checkResult(-3642, 1872);
        nextCycle(3386); checkResult(-3639, 1878);
        nextCycle(3387); checkResult(-3636, 1883);
        nextCycle(3388); checkResult(-3633, 1889);
        nextCycle(3389); checkResult(-3631, 1894);
        nextCycle(3390); checkResult(-3628, 1900);
        nextCycle(3391); checkResult(-3625, 1905);
        nextCycle(3392); checkResult(-3622, 1911);
        nextCycle(3393); checkResult(-3619, 1917);
        nextCycle(3394); checkResult(-3616, 1922);
        nextCycle(3395); checkResult(-3613, 1928);
        nextCycle(3396); checkResult(-3610, 1933);
        nextCycle(3397); checkResult(-3607, 1939);
        nextCycle(3398); checkResult(-3604, 1944);
        nextCycle(3399); checkResult(-3601, 1950);
        nextCycle(3400); checkResult(-3598, 1955);
        nextCycle(3401); checkResult(-3595, 1961);
        nextCycle(3402); checkResult(-3592, 1966);
        nextCycle(3403); checkResult(-3589, 1972);
        nextCycle(3404); checkResult(-3586, 1977);
        nextCycle(3405); checkResult(-3583, 1983);
        nextCycle(3406); checkResult(-3580, 1988);
        nextCycle(3407); checkResult(-3577, 1994);
        nextCycle(3408); checkResult(-3574, 1999);
        nextCycle(3409); checkResult(-3571, 2005);
        nextCycle(3410); checkResult(-3568, 2010);
        nextCycle(3411); checkResult(-3565, 2016);
        nextCycle(3412); checkResult(-3561, 2021);
        nextCycle(3413); checkResult(-3558, 2027);
        nextCycle(3414); checkResult(-3555, 2032);
        nextCycle(3415); checkResult(-3552, 2038);
        nextCycle(3416); checkResult(-3549, 2043);
        nextCycle(3417); checkResult(-3546, 2048);
        nextCycle(3418); checkResult(-3543, 2054);
        nextCycle(3419); checkResult(-3540, 2059);
        nextCycle(3420); checkResult(-3536, 2065);
        nextCycle(3421); checkResult(-3533, 2070);
        nextCycle(3422); checkResult(-3530, 2076);
        nextCycle(3423); checkResult(-3527, 2081);
        nextCycle(3424); checkResult(-3524, 2086);
        nextCycle(3425); checkResult(-3520, 2092);
        nextCycle(3426); checkResult(-3517, 2097);
        nextCycle(3427); checkResult(-3514, 2103);
        nextCycle(3428); checkResult(-3511, 2108);
        nextCycle(3429); checkResult(-3508, 2113);
        nextCycle(3430); checkResult(-3504, 2119);
        nextCycle(3431); checkResult(-3501, 2124);
        nextCycle(3432); checkResult(-3498, 2129);
        nextCycle(3433); checkResult(-3495, 2135);
        nextCycle(3434); checkResult(-3491, 2140);
        nextCycle(3435); checkResult(-3488, 2146);
        nextCycle(3436); checkResult(-3485, 2151);
        nextCycle(3437); checkResult(-3481, 2156);
        nextCycle(3438); checkResult(-3478, 2162);
        nextCycle(3439); checkResult(-3475, 2167);
        nextCycle(3440); checkResult(-3471, 2172);
        nextCycle(3441); checkResult(-3468, 2178);
        nextCycle(3442); checkResult(-3465, 2183);
        nextCycle(3443); checkResult(-3461, 2188);
        nextCycle(3444); checkResult(-3458, 2193);
        nextCycle(3445); checkResult(-3455, 2199);
        nextCycle(3446); checkResult(-3451, 2204);
        nextCycle(3447); checkResult(-3448, 2209);
        nextCycle(3448); checkResult(-3444, 2215);
        nextCycle(3449); checkResult(-3441, 2220);
        nextCycle(3450); checkResult(-3438, 2225);
        nextCycle(3451); checkResult(-3434, 2230);
        nextCycle(3452); checkResult(-3431, 2236);
        nextCycle(3453); checkResult(-3427, 2241);
        nextCycle(3454); checkResult(-3424, 2246);
        nextCycle(3455); checkResult(-3420, 2252);
        nextCycle(3456); checkResult(-3417, 2257);
        nextCycle(3457); checkResult(-3414, 2262);
        nextCycle(3458); checkResult(-3410, 2267);
        nextCycle(3459); checkResult(-3407, 2272);
        nextCycle(3460); checkResult(-3403, 2278);
        nextCycle(3461); checkResult(-3400, 2283);
        nextCycle(3462); checkResult(-3396, 2288);
        nextCycle(3463); checkResult(-3393, 2293);
        nextCycle(3464); checkResult(-3389, 2299);
        nextCycle(3465); checkResult(-3386, 2304);
        nextCycle(3466); checkResult(-3382, 2309);
        nextCycle(3467); checkResult(-3378, 2314);
        nextCycle(3468); checkResult(-3375, 2319);
        nextCycle(3469); checkResult(-3371, 2324);
        nextCycle(3470); checkResult(-3368, 2330);
        nextCycle(3471); checkResult(-3364, 2335);
        nextCycle(3472); checkResult(-3361, 2340);
        nextCycle(3473); checkResult(-3357, 2345);
        nextCycle(3474); checkResult(-3353, 2350);
        nextCycle(3475); checkResult(-3350, 2355);
        nextCycle(3476); checkResult(-3346, 2361);
        nextCycle(3477); checkResult(-3343, 2366);
        nextCycle(3478); checkResult(-3339, 2371);
        nextCycle(3479); checkResult(-3335, 2376);
        nextCycle(3480); checkResult(-3332, 2381);
        nextCycle(3481); checkResult(-3328, 2386);
        nextCycle(3482); checkResult(-3324, 2391);
        nextCycle(3483); checkResult(-3321, 2396);
        nextCycle(3484); checkResult(-3317, 2401);
        nextCycle(3485); checkResult(-3313, 2406);
        nextCycle(3486); checkResult(-3310, 2412);
        nextCycle(3487); checkResult(-3306, 2417);
        nextCycle(3488); checkResult(-3302, 2422);
        nextCycle(3489); checkResult(-3298, 2427);
        nextCycle(3490); checkResult(-3295, 2432);
        nextCycle(3491); checkResult(-3291, 2437);
        nextCycle(3492); checkResult(-3287, 2442);
        nextCycle(3493); checkResult(-3284, 2447);
        nextCycle(3494); checkResult(-3280, 2452);
        nextCycle(3495); checkResult(-3276, 2457);
        nextCycle(3496); checkResult(-3272, 2462);
        nextCycle(3497); checkResult(-3268, 2467);
        nextCycle(3498); checkResult(-3265, 2472);
        nextCycle(3499); checkResult(-3261, 2477);
        nextCycle(3500); checkResult(-3257, 2482);
        nextCycle(3501); checkResult(-3253, 2487);
        nextCycle(3502); checkResult(-3249, 2492);
        nextCycle(3503); checkResult(-3246, 2497);
        nextCycle(3504); checkResult(-3242, 2502);
        nextCycle(3505); checkResult(-3238, 2507);
        nextCycle(3506); checkResult(-3234, 2512);
        nextCycle(3507); checkResult(-3230, 2517);
        nextCycle(3508); checkResult(-3226, 2522);
        nextCycle(3509); checkResult(-3222, 2527);
        nextCycle(3510); checkResult(-3219, 2532);
        nextCycle(3511); checkResult(-3215, 2537);
        nextCycle(3512); checkResult(-3211, 2542);
        nextCycle(3513); checkResult(-3207, 2547);
        nextCycle(3514); checkResult(-3203, 2551);
        nextCycle(3515); checkResult(-3199, 2556);
        nextCycle(3516); checkResult(-3195, 2561);
        nextCycle(3517); checkResult(-3191, 2566);
        nextCycle(3518); checkResult(-3187, 2571);
        nextCycle(3519); checkResult(-3183, 2576);
        nextCycle(3520); checkResult(-3179, 2581);
        nextCycle(3521); checkResult(-3175, 2586);
        nextCycle(3522); checkResult(-3171, 2591);
        nextCycle(3523); checkResult(-3167, 2595);
        nextCycle(3524); checkResult(-3163, 2600);
        nextCycle(3525); checkResult(-3159, 2605);
        nextCycle(3526); checkResult(-3155, 2610);
        nextCycle(3527); checkResult(-3151, 2615);
        nextCycle(3528); checkResult(-3147, 2620);
        nextCycle(3529); checkResult(-3143, 2624);
        nextCycle(3530); checkResult(-3139, 2629);
        nextCycle(3531); checkResult(-3135, 2634);
        nextCycle(3532); checkResult(-3131, 2639);
        nextCycle(3533); checkResult(-3127, 2644);
        nextCycle(3534); checkResult(-3123, 2648);
        nextCycle(3535); checkResult(-3119, 2653);
        nextCycle(3536); checkResult(-3115, 2658);
        nextCycle(3537); checkResult(-3111, 2663);
        nextCycle(3538); checkResult(-3107, 2668);
        nextCycle(3539); checkResult(-3103, 2672);
        nextCycle(3540); checkResult(-3099, 2677);
        nextCycle(3541); checkResult(-3095, 2682);
        nextCycle(3542); checkResult(-3090, 2687);
        nextCycle(3543); checkResult(-3086, 2691);
        nextCycle(3544); checkResult(-3082, 2696);
        nextCycle(3545); checkResult(-3078, 2701);
        nextCycle(3546); checkResult(-3074, 2706);
        nextCycle(3547); checkResult(-3070, 2710);
        nextCycle(3548); checkResult(-3066, 2715);
        nextCycle(3549); checkResult(-3061, 2720);
        nextCycle(3550); checkResult(-3057, 2724);
        nextCycle(3551); checkResult(-3053, 2729);
        nextCycle(3552); checkResult(-3049, 2734);
        nextCycle(3553); checkResult(-3045, 2738);
        nextCycle(3554); checkResult(-3041, 2743);
        nextCycle(3555); checkResult(-3036, 2748);
        nextCycle(3556); checkResult(-3032, 2752);
        nextCycle(3557); checkResult(-3028, 2757);
        nextCycle(3558); checkResult(-3024, 2762);
        nextCycle(3559); checkResult(-3019, 2766);
        nextCycle(3560); checkResult(-3015, 2771);
        nextCycle(3561); checkResult(-3011, 2776);
        nextCycle(3562); checkResult(-3007, 2780);
        nextCycle(3563); checkResult(-3002, 2785);
        nextCycle(3564); checkResult(-2998, 2789);
        nextCycle(3565); checkResult(-2994, 2794);
        nextCycle(3566); checkResult(-2990, 2799);
        nextCycle(3567); checkResult(-2985, 2803);
        nextCycle(3568); checkResult(-2981, 2808);
        nextCycle(3569); checkResult(-2977, 2812);
        nextCycle(3570); checkResult(-2972, 2817);
        nextCycle(3571); checkResult(-2968, 2821);
        nextCycle(3572); checkResult(-2964, 2826);
        nextCycle(3573); checkResult(-2959, 2830);
        nextCycle(3574); checkResult(-2955, 2835);
        nextCycle(3575); checkResult(-2951, 2840);
        nextCycle(3576); checkResult(-2946, 2844);
        nextCycle(3577); checkResult(-2942, 2849);
        nextCycle(3578); checkResult(-2937, 2853);
        nextCycle(3579); checkResult(-2933, 2858);
        nextCycle(3580); checkResult(-2929, 2862);
        nextCycle(3581); checkResult(-2924, 2867);
        nextCycle(3582); checkResult(-2920, 2871);
        nextCycle(3583); checkResult(-2916, 2876);
        nextCycle(3584); checkResult(-2911, 2880);
        nextCycle(3585); checkResult(-2907, 2884);
        nextCycle(3586); checkResult(-2902, 2889);
        nextCycle(3587); checkResult(-2898, 2893);
        nextCycle(3588); checkResult(-2893, 2898);
        nextCycle(3589); checkResult(-2889, 2902);
        nextCycle(3590); checkResult(-2884, 2907);
        nextCycle(3591); checkResult(-2880, 2911);
        nextCycle(3592); checkResult(-2876, 2916);
        nextCycle(3593); checkResult(-2871, 2920);
        nextCycle(3594); checkResult(-2867, 2924);
        nextCycle(3595); checkResult(-2862, 2929);
        nextCycle(3596); checkResult(-2858, 2933);
        nextCycle(3597); checkResult(-2853, 2937);
        nextCycle(3598); checkResult(-2849, 2942);
        nextCycle(3599); checkResult(-2844, 2946);
        nextCycle(3600); checkResult(-2840, 2951);
        nextCycle(3601); checkResult(-2835, 2955);
        nextCycle(3602); checkResult(-2830, 2959);
        nextCycle(3603); checkResult(-2826, 2964);
        nextCycle(3604); checkResult(-2821, 2968);
        nextCycle(3605); checkResult(-2817, 2972);
        nextCycle(3606); checkResult(-2812, 2977);
        nextCycle(3607); checkResult(-2808, 2981);
        nextCycle(3608); checkResult(-2803, 2985);
        nextCycle(3609); checkResult(-2799, 2990);
        nextCycle(3610); checkResult(-2794, 2994);
        nextCycle(3611); checkResult(-2789, 2998);
        nextCycle(3612); checkResult(-2785, 3002);
        nextCycle(3613); checkResult(-2780, 3007);
        nextCycle(3614); checkResult(-2776, 3011);
        nextCycle(3615); checkResult(-2771, 3015);
        nextCycle(3616); checkResult(-2766, 3019);
        nextCycle(3617); checkResult(-2762, 3024);
        nextCycle(3618); checkResult(-2757, 3028);
        nextCycle(3619); checkResult(-2752, 3032);
        nextCycle(3620); checkResult(-2748, 3036);
        nextCycle(3621); checkResult(-2743, 3041);
        nextCycle(3622); checkResult(-2738, 3045);
        nextCycle(3623); checkResult(-2734, 3049);
        nextCycle(3624); checkResult(-2729, 3053);
        nextCycle(3625); checkResult(-2724, 3057);
        nextCycle(3626); checkResult(-2720, 3061);
        nextCycle(3627); checkResult(-2715, 3066);
        nextCycle(3628); checkResult(-2710, 3070);
        nextCycle(3629); checkResult(-2706, 3074);
        nextCycle(3630); checkResult(-2701, 3078);
        nextCycle(3631); checkResult(-2696, 3082);
        nextCycle(3632); checkResult(-2691, 3086);
        nextCycle(3633); checkResult(-2687, 3090);
        nextCycle(3634); checkResult(-2682, 3095);
        nextCycle(3635); checkResult(-2677, 3099);
        nextCycle(3636); checkResult(-2672, 3103);
        nextCycle(3637); checkResult(-2668, 3107);
        nextCycle(3638); checkResult(-2663, 3111);
        nextCycle(3639); checkResult(-2658, 3115);
        nextCycle(3640); checkResult(-2653, 3119);
        nextCycle(3641); checkResult(-2648, 3123);
        nextCycle(3642); checkResult(-2644, 3127);
        nextCycle(3643); checkResult(-2639, 3131);
        nextCycle(3644); checkResult(-2634, 3135);
        nextCycle(3645); checkResult(-2629, 3139);
        nextCycle(3646); checkResult(-2624, 3143);
        nextCycle(3647); checkResult(-2620, 3147);
        nextCycle(3648); checkResult(-2615, 3151);
        nextCycle(3649); checkResult(-2610, 3155);
        nextCycle(3650); checkResult(-2605, 3159);
        nextCycle(3651); checkResult(-2600, 3163);
        nextCycle(3652); checkResult(-2595, 3167);
        nextCycle(3653); checkResult(-2591, 3171);
        nextCycle(3654); checkResult(-2586, 3175);
        nextCycle(3655); checkResult(-2581, 3179);
        nextCycle(3656); checkResult(-2576, 3183);
        nextCycle(3657); checkResult(-2571, 3187);
        nextCycle(3658); checkResult(-2566, 3191);
        nextCycle(3659); checkResult(-2561, 3195);
        nextCycle(3660); checkResult(-2556, 3199);
        nextCycle(3661); checkResult(-2551, 3203);
        nextCycle(3662); checkResult(-2547, 3207);
        nextCycle(3663); checkResult(-2542, 3211);
        nextCycle(3664); checkResult(-2537, 3215);
        nextCycle(3665); checkResult(-2532, 3219);
        nextCycle(3666); checkResult(-2527, 3222);
        nextCycle(3667); checkResult(-2522, 3226);
        nextCycle(3668); checkResult(-2517, 3230);
        nextCycle(3669); checkResult(-2512, 3234);
        nextCycle(3670); checkResult(-2507, 3238);
        nextCycle(3671); checkResult(-2502, 3242);
        nextCycle(3672); checkResult(-2497, 3246);
        nextCycle(3673); checkResult(-2492, 3249);
        nextCycle(3674); checkResult(-2487, 3253);
        nextCycle(3675); checkResult(-2482, 3257);
        nextCycle(3676); checkResult(-2477, 3261);
        nextCycle(3677); checkResult(-2472, 3265);
        nextCycle(3678); checkResult(-2467, 3268);
        nextCycle(3679); checkResult(-2462, 3272);
        nextCycle(3680); checkResult(-2457, 3276);
        nextCycle(3681); checkResult(-2452, 3280);
        nextCycle(3682); checkResult(-2447, 3284);
        nextCycle(3683); checkResult(-2442, 3287);
        nextCycle(3684); checkResult(-2437, 3291);
        nextCycle(3685); checkResult(-2432, 3295);
        nextCycle(3686); checkResult(-2427, 3298);
        nextCycle(3687); checkResult(-2422, 3302);
        nextCycle(3688); checkResult(-2417, 3306);
        nextCycle(3689); checkResult(-2412, 3310);
        nextCycle(3690); checkResult(-2406, 3313);
        nextCycle(3691); checkResult(-2401, 3317);
        nextCycle(3692); checkResult(-2396, 3321);
        nextCycle(3693); checkResult(-2391, 3324);
        nextCycle(3694); checkResult(-2386, 3328);
        nextCycle(3695); checkResult(-2381, 3332);
        nextCycle(3696); checkResult(-2376, 3335);
        nextCycle(3697); checkResult(-2371, 3339);
        nextCycle(3698); checkResult(-2366, 3343);
        nextCycle(3699); checkResult(-2361, 3346);
        nextCycle(3700); checkResult(-2355, 3350);
        nextCycle(3701); checkResult(-2350, 3353);
        nextCycle(3702); checkResult(-2345, 3357);
        nextCycle(3703); checkResult(-2340, 3361);
        nextCycle(3704); checkResult(-2335, 3364);
        nextCycle(3705); checkResult(-2330, 3368);
        nextCycle(3706); checkResult(-2324, 3371);
        nextCycle(3707); checkResult(-2319, 3375);
        nextCycle(3708); checkResult(-2314, 3378);
        nextCycle(3709); checkResult(-2309, 3382);
        nextCycle(3710); checkResult(-2304, 3386);
        nextCycle(3711); checkResult(-2299, 3389);
        nextCycle(3712); checkResult(-2293, 3393);
        nextCycle(3713); checkResult(-2288, 3396);
        nextCycle(3714); checkResult(-2283, 3400);
        nextCycle(3715); checkResult(-2278, 3403);
        nextCycle(3716); checkResult(-2272, 3407);
        nextCycle(3717); checkResult(-2267, 3410);
        nextCycle(3718); checkResult(-2262, 3414);
        nextCycle(3719); checkResult(-2257, 3417);
        nextCycle(3720); checkResult(-2252, 3420);
        nextCycle(3721); checkResult(-2246, 3424);
        nextCycle(3722); checkResult(-2241, 3427);
        nextCycle(3723); checkResult(-2236, 3431);
        nextCycle(3724); checkResult(-2230, 3434);
        nextCycle(3725); checkResult(-2225, 3438);
        nextCycle(3726); checkResult(-2220, 3441);
        nextCycle(3727); checkResult(-2215, 3444);
        nextCycle(3728); checkResult(-2209, 3448);
        nextCycle(3729); checkResult(-2204, 3451);
        nextCycle(3730); checkResult(-2199, 3455);
        nextCycle(3731); checkResult(-2193, 3458);
        nextCycle(3732); checkResult(-2188, 3461);
        nextCycle(3733); checkResult(-2183, 3465);
        nextCycle(3734); checkResult(-2178, 3468);
        nextCycle(3735); checkResult(-2172, 3471);
        nextCycle(3736); checkResult(-2167, 3475);
        nextCycle(3737); checkResult(-2162, 3478);
        nextCycle(3738); checkResult(-2156, 3481);
        nextCycle(3739); checkResult(-2151, 3485);
        nextCycle(3740); checkResult(-2146, 3488);
        nextCycle(3741); checkResult(-2140, 3491);
        nextCycle(3742); checkResult(-2135, 3495);
        nextCycle(3743); checkResult(-2129, 3498);
        nextCycle(3744); checkResult(-2124, 3501);
        nextCycle(3745); checkResult(-2119, 3504);
        nextCycle(3746); checkResult(-2113, 3508);
        nextCycle(3747); checkResult(-2108, 3511);
        nextCycle(3748); checkResult(-2103, 3514);
        nextCycle(3749); checkResult(-2097, 3517);
        nextCycle(3750); checkResult(-2092, 3520);
        nextCycle(3751); checkResult(-2086, 3524);
        nextCycle(3752); checkResult(-2081, 3527);
        nextCycle(3753); checkResult(-2076, 3530);
        nextCycle(3754); checkResult(-2070, 3533);
        nextCycle(3755); checkResult(-2065, 3536);
        nextCycle(3756); checkResult(-2059, 3540);
        nextCycle(3757); checkResult(-2054, 3543);
        nextCycle(3758); checkResult(-2048, 3546);
        nextCycle(3759); checkResult(-2043, 3549);
        nextCycle(3760); checkResult(-2038, 3552);
        nextCycle(3761); checkResult(-2032, 3555);
        nextCycle(3762); checkResult(-2027, 3558);
        nextCycle(3763); checkResult(-2021, 3561);
        nextCycle(3764); checkResult(-2016, 3565);
        nextCycle(3765); checkResult(-2010, 3568);
        nextCycle(3766); checkResult(-2005, 3571);
        nextCycle(3767); checkResult(-1999, 3574);
        nextCycle(3768); checkResult(-1994, 3577);
        nextCycle(3769); checkResult(-1988, 3580);
        nextCycle(3770); checkResult(-1983, 3583);
        nextCycle(3771); checkResult(-1977, 3586);
        nextCycle(3772); checkResult(-1972, 3589);
        nextCycle(3773); checkResult(-1966, 3592);
        nextCycle(3774); checkResult(-1961, 3595);
        nextCycle(3775); checkResult(-1955, 3598);
        nextCycle(3776); checkResult(-1950, 3601);
        nextCycle(3777); checkResult(-1944, 3604);
        nextCycle(3778); checkResult(-1939, 3607);
        nextCycle(3779); checkResult(-1933, 3610);
        nextCycle(3780); checkResult(-1928, 3613);
        nextCycle(3781); checkResult(-1922, 3616);
        nextCycle(3782); checkResult(-1917, 3619);
        nextCycle(3783); checkResult(-1911, 3622);
        nextCycle(3784); checkResult(-1905, 3625);
        nextCycle(3785); checkResult(-1900, 3628);
        nextCycle(3786); checkResult(-1894, 3631);
        nextCycle(3787); checkResult(-1889, 3633);
        nextCycle(3788); checkResult(-1883, 3636);
        nextCycle(3789); checkResult(-1878, 3639);
        nextCycle(3790); checkResult(-1872, 3642);
        nextCycle(3791); checkResult(-1866, 3645);
        nextCycle(3792); checkResult(-1861, 3648);
        nextCycle(3793); checkResult(-1855, 3651);
        nextCycle(3794); checkResult(-1850, 3654);
        nextCycle(3795); checkResult(-1844, 3656);
        nextCycle(3796); checkResult(-1838, 3659);
        nextCycle(3797); checkResult(-1833, 3662);
        nextCycle(3798); checkResult(-1827, 3665);
        nextCycle(3799); checkResult(-1821, 3668);
        nextCycle(3800); checkResult(-1816, 3670);
        nextCycle(3801); checkResult(-1810, 3673);
        nextCycle(3802); checkResult(-1805, 3676);
        nextCycle(3803); checkResult(-1799, 3679);
        nextCycle(3804); checkResult(-1793, 3681);
        nextCycle(3805); checkResult(-1788, 3684);
        nextCycle(3806); checkResult(-1782, 3687);
        nextCycle(3807); checkResult(-1776, 3690);
        nextCycle(3808); checkResult(-1771, 3692);
        nextCycle(3809); checkResult(-1765, 3695);
        nextCycle(3810); checkResult(-1759, 3698);
        nextCycle(3811); checkResult(-1754, 3700);
        nextCycle(3812); checkResult(-1748, 3703);
        nextCycle(3813); checkResult(-1742, 3706);
        nextCycle(3814); checkResult(-1737, 3709);
        nextCycle(3815); checkResult(-1731, 3711);
        nextCycle(3816); checkResult(-1725, 3714);
        nextCycle(3817); checkResult(-1720, 3716);
        nextCycle(3818); checkResult(-1714, 3719);
        nextCycle(3819); checkResult(-1708, 3722);
        nextCycle(3820); checkResult(-1702, 3724);
        nextCycle(3821); checkResult(-1697, 3727);
        nextCycle(3822); checkResult(-1691, 3730);
        nextCycle(3823); checkResult(-1685, 3732);
        nextCycle(3824); checkResult(-1680, 3735);
        nextCycle(3825); checkResult(-1674, 3737);
        nextCycle(3826); checkResult(-1668, 3740);
        nextCycle(3827); checkResult(-1662, 3742);
        nextCycle(3828); checkResult(-1657, 3745);
        nextCycle(3829); checkResult(-1651, 3747);
        nextCycle(3830); checkResult(-1645, 3750);
        nextCycle(3831); checkResult(-1639, 3753);
        nextCycle(3832); checkResult(-1634, 3755);
        nextCycle(3833); checkResult(-1628, 3758);
        nextCycle(3834); checkResult(-1622, 3760);
        nextCycle(3835); checkResult(-1616, 3763);
        nextCycle(3836); checkResult(-1611, 3765);
        nextCycle(3837); checkResult(-1605, 3767);
        nextCycle(3838); checkResult(-1599, 3770);
        nextCycle(3839); checkResult(-1593, 3772);
        nextCycle(3840); checkResult(-1587, 3775);
        nextCycle(3841); checkResult(-1582, 3777);
        nextCycle(3842); checkResult(-1576, 3780);
        nextCycle(3843); checkResult(-1570, 3782);
        nextCycle(3844); checkResult(-1564, 3784);
        nextCycle(3845); checkResult(-1558, 3787);
        nextCycle(3846); checkResult(-1553, 3789);
        nextCycle(3847); checkResult(-1547, 3792);
        nextCycle(3848); checkResult(-1541, 3794);
        nextCycle(3849); checkResult(-1535, 3796);
        nextCycle(3850); checkResult(-1529, 3799);
        nextCycle(3851); checkResult(-1523, 3801);
        nextCycle(3852); checkResult(-1518, 3803);
        nextCycle(3853); checkResult(-1512, 3806);
        nextCycle(3854); checkResult(-1506, 3808);
        nextCycle(3855); checkResult(-1500, 3810);
        nextCycle(3856); checkResult(-1494, 3813);
        nextCycle(3857); checkResult(-1488, 3815);
        nextCycle(3858); checkResult(-1483, 3817);
        nextCycle(3859); checkResult(-1477, 3819);
        nextCycle(3860); checkResult(-1471, 3822);
        nextCycle(3861); checkResult(-1465, 3824);
        nextCycle(3862); checkResult(-1459, 3826);
        nextCycle(3863); checkResult(-1453, 3828);
        nextCycle(3864); checkResult(-1447, 3831);
        nextCycle(3865); checkResult(-1441, 3833);
        nextCycle(3866); checkResult(-1436, 3835);
        nextCycle(3867); checkResult(-1430, 3837);
        nextCycle(3868); checkResult(-1424, 3839);
        nextCycle(3869); checkResult(-1418, 3842);
        nextCycle(3870); checkResult(-1412, 3844);
        nextCycle(3871); checkResult(-1406, 3846);
        nextCycle(3872); checkResult(-1400, 3848);
        nextCycle(3873); checkResult(-1394, 3850);
        nextCycle(3874); checkResult(-1388, 3852);
        nextCycle(3875); checkResult(-1383, 3855);
        nextCycle(3876); checkResult(-1377, 3857);
        nextCycle(3877); checkResult(-1371, 3859);
        nextCycle(3878); checkResult(-1365, 3861);
        nextCycle(3879); checkResult(-1359, 3863);
        nextCycle(3880); checkResult(-1353, 3865);
        nextCycle(3881); checkResult(-1347, 3867);
        nextCycle(3882); checkResult(-1341, 3869);
        nextCycle(3883); checkResult(-1335, 3871);
        nextCycle(3884); checkResult(-1329, 3873);
        nextCycle(3885); checkResult(-1323, 3875);
        nextCycle(3886); checkResult(-1317, 3877);
        nextCycle(3887); checkResult(-1311, 3879);
        nextCycle(3888); checkResult(-1305, 3881);
        nextCycle(3889); checkResult(-1299, 3883);
        nextCycle(3890); checkResult(-1293, 3885);
        nextCycle(3891); checkResult(-1288, 3887);
        nextCycle(3892); checkResult(-1282, 3889);
        nextCycle(3893); checkResult(-1276, 3891);
        nextCycle(3894); checkResult(-1270, 3893);
        nextCycle(3895); checkResult(-1264, 3895);
        nextCycle(3896); checkResult(-1258, 3897);
        nextCycle(3897); checkResult(-1252, 3899);
        nextCycle(3898); checkResult(-1246, 3901);
        nextCycle(3899); checkResult(-1240, 3903);
        nextCycle(3900); checkResult(-1234, 3905);
        nextCycle(3901); checkResult(-1228, 3907);
        nextCycle(3902); checkResult(-1222, 3909);
        nextCycle(3903); checkResult(-1216, 3910);
        nextCycle(3904); checkResult(-1210, 3912);
        nextCycle(3905); checkResult(-1204, 3914);
        nextCycle(3906); checkResult(-1198, 3916);
        nextCycle(3907); checkResult(-1192, 3918);
        nextCycle(3908); checkResult(-1186, 3920);
        nextCycle(3909); checkResult(-1180, 3921);
        nextCycle(3910); checkResult(-1174, 3923);
        nextCycle(3911); checkResult(-1168, 3925);
        nextCycle(3912); checkResult(-1162, 3927);
        nextCycle(3913); checkResult(-1156, 3929);
        nextCycle(3914); checkResult(-1150, 3930);
        nextCycle(3915); checkResult(-1144, 3932);
        nextCycle(3916); checkResult(-1138, 3934);
        nextCycle(3917); checkResult(-1131, 3936);
        nextCycle(3918); checkResult(-1125, 3937);
        nextCycle(3919); checkResult(-1119, 3939);
        nextCycle(3920); checkResult(-1113, 3941);
        nextCycle(3921); checkResult(-1107, 3942);
        nextCycle(3922); checkResult(-1101, 3944);
        nextCycle(3923); checkResult(-1095, 3946);
        nextCycle(3924); checkResult(-1089, 3947);
        nextCycle(3925); checkResult(-1083, 3949);
        nextCycle(3926); checkResult(-1077, 3951);
        nextCycle(3927); checkResult(-1071, 3952);
        nextCycle(3928); checkResult(-1065, 3954);
        nextCycle(3929); checkResult(-1059, 3956);
        nextCycle(3930); checkResult(-1053, 3957);
        nextCycle(3931); checkResult(-1047, 3959);
        nextCycle(3932); checkResult(-1041, 3961);
        nextCycle(3933); checkResult(-1035, 3962);
        nextCycle(3934); checkResult(-1028, 3964);
        nextCycle(3935); checkResult(-1022, 3965);
        nextCycle(3936); checkResult(-1016, 3967);
        nextCycle(3937); checkResult(-1010, 3968);
        nextCycle(3938); checkResult(-1004, 3970);
        nextCycle(3939); checkResult(-998, 3972);
        nextCycle(3940); checkResult(-992, 3973);
        nextCycle(3941); checkResult(-986, 3975);
        nextCycle(3942); checkResult(-980, 3976);
        nextCycle(3943); checkResult(-974, 3978);
        nextCycle(3944); checkResult(-968, 3979);
        nextCycle(3945); checkResult(-961, 3981);
        nextCycle(3946); checkResult(-955, 3982);
        nextCycle(3947); checkResult(-949, 3983);
        nextCycle(3948); checkResult(-943, 3985);
        nextCycle(3949); checkResult(-937, 3986);
        nextCycle(3950); checkResult(-931, 3988);
        nextCycle(3951); checkResult(-925, 3989);
        nextCycle(3952); checkResult(-919, 3991);
        nextCycle(3953); checkResult(-913, 3992);
        nextCycle(3954); checkResult(-906, 3993);
        nextCycle(3955); checkResult(-900, 3995);
        nextCycle(3956); checkResult(-894, 3996);
        nextCycle(3957); checkResult(-888, 3998);
        nextCycle(3958); checkResult(-882, 3999);
        nextCycle(3959); checkResult(-876, 4000);
        nextCycle(3960); checkResult(-870, 4002);
        nextCycle(3961); checkResult(-863, 4003);
        nextCycle(3962); checkResult(-857, 4004);
        nextCycle(3963); checkResult(-851, 4006);
        nextCycle(3964); checkResult(-845, 4007);
        nextCycle(3965); checkResult(-839, 4008);
        nextCycle(3966); checkResult(-833, 4009);
        nextCycle(3967); checkResult(-827, 4011);
        nextCycle(3968); checkResult(-820, 4012);
        nextCycle(3969); checkResult(-814, 4013);
        nextCycle(3970); checkResult(-808, 4014);
        nextCycle(3971); checkResult(-802, 4016);
        nextCycle(3972); checkResult(-796, 4017);
        nextCycle(3973); checkResult(-790, 4018);
        nextCycle(3974); checkResult(-783, 4019);
        nextCycle(3975); checkResult(-777, 4021);
        nextCycle(3976); checkResult(-771, 4022);
        nextCycle(3977); checkResult(-765, 4023);
        nextCycle(3978); checkResult(-759, 4024);
        nextCycle(3979); checkResult(-753, 4025);
        nextCycle(3980); checkResult(-746, 4026);
        nextCycle(3981); checkResult(-740, 4028);
        nextCycle(3982); checkResult(-734, 4029);
        nextCycle(3983); checkResult(-728, 4030);
        nextCycle(3984); checkResult(-722, 4031);
        nextCycle(3985); checkResult(-716, 4032);
        nextCycle(3986); checkResult(-709, 4033);
        nextCycle(3987); checkResult(-703, 4034);
        nextCycle(3988); checkResult(-697, 4035);
        nextCycle(3989); checkResult(-691, 4036);
        nextCycle(3990); checkResult(-685, 4037);
        nextCycle(3991); checkResult(-678, 4038);
        nextCycle(3992); checkResult(-672, 4039);
        nextCycle(3993); checkResult(-666, 4040);
        nextCycle(3994); checkResult(-660, 4041);
        nextCycle(3995); checkResult(-654, 4042);
        nextCycle(3996); checkResult(-647, 4043);
        nextCycle(3997); checkResult(-641, 4044);
        nextCycle(3998); checkResult(-635, 4045);
        nextCycle(3999); checkResult(-629, 4046);
        nextCycle(4000); checkResult(-623, 4047);
        nextCycle(4001); checkResult(-616, 4048);
        nextCycle(4002); checkResult(-610, 4049);
        nextCycle(4003); checkResult(-604, 4050);
        nextCycle(4004); checkResult(-598, 4051);
        nextCycle(4005); checkResult(-592, 4052);
        nextCycle(4006); checkResult(-585, 4053);
        nextCycle(4007); checkResult(-579, 4054);
        nextCycle(4008); checkResult(-573, 4055);
        nextCycle(4009); checkResult(-567, 4056);
        nextCycle(4010); checkResult(-560, 4056);
        nextCycle(4011); checkResult(-554, 4057);
        nextCycle(4012); checkResult(-548, 4058);
        nextCycle(4013); checkResult(-542, 4059);
        nextCycle(4014); checkResult(-536, 4060);
        nextCycle(4015); checkResult(-529, 4061);
        nextCycle(4016); checkResult(-523, 4061);
        nextCycle(4017); checkResult(-517, 4062);
        nextCycle(4018); checkResult(-511, 4063);
        nextCycle(4019); checkResult(-504, 4064);
        nextCycle(4020); checkResult(-498, 4065);
        nextCycle(4021); checkResult(-492, 4065);
        nextCycle(4022); checkResult(-486, 4066);
        nextCycle(4023); checkResult(-479, 4067);
        nextCycle(4024); checkResult(-473, 4068);
        nextCycle(4025); checkResult(-467, 4068);
        nextCycle(4026); checkResult(-461, 4069);
        nextCycle(4027); checkResult(-454, 4070);
        nextCycle(4028); checkResult(-448, 4070);
        nextCycle(4029); checkResult(-442, 4071);
        nextCycle(4030); checkResult(-436, 4072);
        nextCycle(4031); checkResult(-430, 4072);
        nextCycle(4032); checkResult(-423, 4073);
        nextCycle(4033); checkResult(-417, 4074);
        nextCycle(4034); checkResult(-411, 4074);
        nextCycle(4035); checkResult(-405, 4075);
        nextCycle(4036); checkResult(-398, 4076);
        nextCycle(4037); checkResult(-392, 4076);
        nextCycle(4038); checkResult(-386, 4077);
        nextCycle(4039); checkResult(-379, 4077);
        nextCycle(4040); checkResult(-373, 4078);
        nextCycle(4041); checkResult(-367, 4079);
        nextCycle(4042); checkResult(-361, 4079);
        nextCycle(4043); checkResult(-354, 4080);
        nextCycle(4044); checkResult(-348, 4080);
        nextCycle(4045); checkResult(-342, 4081);
        nextCycle(4046); checkResult(-336, 4081);
        nextCycle(4047); checkResult(-329, 4082);
        nextCycle(4048); checkResult(-323, 4082);
        nextCycle(4049); checkResult(-317, 4083);
        nextCycle(4050); checkResult(-311, 4083);
        nextCycle(4051); checkResult(-304, 4084);
        nextCycle(4052); checkResult(-298, 4084);
        nextCycle(4053); checkResult(-292, 4085);
        nextCycle(4054); checkResult(-286, 4085);
        nextCycle(4055); checkResult(-279, 4085);
        nextCycle(4056); checkResult(-273, 4086);
        nextCycle(4057); checkResult(-267, 4086);
        nextCycle(4058); checkResult(-261, 4087);
        nextCycle(4059); checkResult(-254, 4087);
        nextCycle(4060); checkResult(-248, 4087);
        nextCycle(4061); checkResult(-242, 4088);
        nextCycle(4062); checkResult(-235, 4088);
        nextCycle(4063); checkResult(-229, 4089);
        nextCycle(4064); checkResult(-223, 4089);
        nextCycle(4065); checkResult(-217, 4089);
        nextCycle(4066); checkResult(-210, 4090);
        nextCycle(4067); checkResult(-204, 4090);
        nextCycle(4068); checkResult(-198, 4090);
        nextCycle(4069); checkResult(-192, 4091);
        nextCycle(4070); checkResult(-185, 4091);
        nextCycle(4071); checkResult(-179, 4091);
        nextCycle(4072); checkResult(-173, 4091);
        nextCycle(4073); checkResult(-166, 4092);
        nextCycle(4074); checkResult(-160, 4092);
        nextCycle(4075); checkResult(-154, 4092);
        nextCycle(4076); checkResult(-148, 4092);
        nextCycle(4077); checkResult(-141, 4093);
        nextCycle(4078); checkResult(-135, 4093);
        nextCycle(4079); checkResult(-129, 4093);
        nextCycle(4080); checkResult(-122, 4093);
        nextCycle(4081); checkResult(-116, 4093);
        nextCycle(4082); checkResult(-110, 4094);
        nextCycle(4083); checkResult(-104, 4094);
        nextCycle(4084); checkResult(-97, 4094);
        nextCycle(4085); checkResult(-91, 4094);
        nextCycle(4086); checkResult(-85, 4094);
        nextCycle(4087); checkResult(-79, 4094);
        nextCycle(4088); checkResult(-72, 4094);
        nextCycle(4089); checkResult(-66, 4094);
        nextCycle(4090); checkResult(-60, 4095);
        nextCycle(4091); checkResult(-53, 4095);
        nextCycle(4092); checkResult(-47, 4095);
        nextCycle(4093); checkResult(-41, 4095);
        nextCycle(4094); checkResult(-35, 4095);
        nextCycle(4095); checkResult(-28, 4095);
        nextCycle(0); checkResult(-22, 4095);
        nextCycle(1); checkResult(-16, 4095);
        nextCycle(2); checkResult(-9, 4095);
        nextCycle(3); checkResult(-3, 4095);
        nextCycle(4); checkResult(3, 4095);
        nextCycle(5); checkResult(9, 4095);
        nextCycle(6); checkResult(16, 4095);
        nextCycle(7); checkResult(22, 4095);
        $display("Test passed");
        $finish();
    end
    
    endmodule
    
