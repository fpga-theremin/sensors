* ADCMP601 SPICE Macro-model
*   06/26 Draft
* LPS APPS Engineering
*
* This is not the final version of ADCMP601 Spice model
*
* This model was created based on the HSPICE version of ADCMP601 by JAV on 6/25/2018
* The ADCMP601 HSPICE model was modified so it can be used in LT SPICE simulator
* This Spice model still needs to be tested to gurantee that it matches the HSPICE version
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | latch/hysteresis
*                | | | positive supply
*                | | | | negative supply
*                | | | | | output pin
*                | | | | | |
*                | | | | | |
*                | | | | | |
.SUBCKT ADCMP601 3 4 5 6 2 1
c0 17 0 5e-13
c1 19 0 2e-13
c2 3 0 2e-13
c3 4 0 2e-13
dp 2 6 DESD
e0 18 0 VALUE = {LIMIT (4*V(17,0),0.3,-0.3)}
e1 20 0 VALUE = {LIMIT (1*V(19,0),0.3,-0.3)}
g0 6 2 0 22 1
io 12 13 dc 1e-06
iq 22 0 dc 0.002422
r0 17 0 700
r1 18 19 1000
r2 3 13 100
r3 4 11 100
r4 21 0 50
rd 3 4 1e7
rp 6 2 1e5
rt 22 0 1 tc=0.0005
t0 20 0 21 0 z0=50 td=1.370e-9
vo 11 12 dc 0.001
x1 4 2 6 ADCMP601_ESD
x2 3 2 6 ADCMP601_ESD
x3 5 2 6 ADCMP601_ESD
x4 1 2 6 ADCMP601_ESD
xb 12 13 14 15 16 2 6 ADCMP601_BIAS
xh 17 2 5 6 ADCMP601_HYST
xi 12 13 14 15 16 17 2 6 ADCMP601_INPUT
xo 1 2 21 6 ADCMP601_OUTPUT
xv 12 13 17 2 6 ADCMP601_DVOS
.ENDS ADCMP601

*
* Bias Current Generator
*
.SUBCKT ADCMP601_BIAS 12 13 14 15 16 2 6
d0 201 202 DSIM1
d1 201 203 DSIM1
d2 205 206 DSIM1
d3 202 204 DSIM1
d4 203 204 DSIM1
d5 207 208 DSIM1
e0 203 0 13 0 1
e1 202 0 12 0 1
e2 205 0 201 0 1
e3 208 0 204 0 1
e4 210 0 VALUE = {LIMIT (1*V(6,209),1.6,0.6)}
e5 219 0 VALUE = {LIMIT (5*V(211,207),1,0)}
g0 2 6 VALUE = {LIMIT (0.0015*V(212,213),0.003,0)}
g1 15 0 VALUE = {LIMIT (0.001*V(212,213),0.002,0)}
g2 16 0 VALUE = {LIMIT (0.001*V(214,215),0.002,0)}
g3 16 0 VALUE = {LIMIT (-0.001*V(214,216),0,-0.0002)}
g4 0 14 VALUE = {LIMIT (0.002*V(217,218),1e-4,0)}
*I=(0+0*V(219,220))+(0+0.2*V(217,218))
g5 6 2 VALUE = {LIMIT (0.002*V(217,218),5e-05,0)}
i0 0 201 dc 0.001
i1 204 0 dc 0.001
i5 206 0 dc 0.001
i6 0 207 dc 0.001
r0 206 218 1
r1 220 0 1
v0 209 0 dc 1.9
v1 211 0 dc 1.6
v2 217 210 dc 0.2
v3 212 207 dc 0.025
v4 213 0 dc 1.6
v5 214 207 dc 0.025
v6 215 0 dc 0.6
v7 216 0 dc 1.7
.ENDS

*
* CMRR and PSRR Offset Generator
*
.SUBCKT ADCMP601_DVOS 12 13 17 2 6
e0 302 0 13 0 1
e1 304 0 12 0 1
g0 17 0 VALUE = {LIMIT (1.71e-06 - 3.3e-07*V(303,0),3e-06,-1e-06)}
*I = 1.71e-06 -3.3e-07*V(303,0)
g1 17 0 VALUE = {LIMIT (6.667e-07*V(6,301),2e-06,0)}
r0 302 303 1000
r1 303 304 1000
v0 301 2 dc 2.5
.ENDS

*
* ESD Diodes
*
.SUBCKT ADCMP601_ESD 601 602 606
d0 601 606 DESD
d1 602 601 DESD
.ENDS

*
* Hysteresis and Latch Function
*
.SUBCKT ADCMP601_HYST 17 2 5 6
c0 410 409 3.4e-11
c1 401 0 1e-12
d0 0 404 DSIM1
d1 401 5 DSIM3
e0 402 405 405 403 1
e1 412 0 VALUE = {LIMIT (20*V(17,0),0.3,-0.3)}
f1 6 0 VALUE = {LIMIT (7*I(v1),0.0007,0)}
f2 0 2 VALUE = {LIMIT (8*I(v2),0.0008,0)}
g0 408 17 VALUE = {LIMIT (0.01*V(410,409),0.0003,-0.0003)}
g1 411 0 VALUE = {LIMIT (0.01*V(414,0),3e-4,0)}
h0 413 0 VALUE = {LIMIT (1000*I(v0),0.030,0)}
i2 403 0 dc 0.00125
i3 5 0 dc 1.25e-06
i5 0 405 dc 1e-06
q0 410 0 411 0 NPN_IN1
q1 409 412 411 0 NPN_IN1
r0 403 404 1000
r1 402 401 7500
r3 408 410 100
r4 408 409 100
r5 414 0 50
t0 413 0 414 0 z0=50 td=7e-10
v0 406 405 0
v1 407 406 0
v2 0 407 0
v4 408 0 dc 1
.ENDS

*
* Input Stage
*
.SUBCKT ADCMP601_INPUT 12 13 14 15 16 17 2 6
e0 101 0 0 2 -1
e1 102 0 0 6 -1
g0 102 17 poly(3) 108 107 106 105 104 103 0 0.01 0.01 0.01
q0 103 13 14 0 PNP_IN1
q1 104 12 14 0 PNP_IN1
q2 105 13 15 0 NPN_IN1
q3 106 12 15 0 NPN_IN1
q4 107 13 16 0 NPN_IN2
q5 108 12 16 0 NPN_IN2
r0 101 103 200
r1 101 104 200
r2 102 105 90
r3 102 106 90
r4 102 107 80
r5 102 108 80
.ENDS

*
* Output Stage
*
.SUBCKT ADCMP601_OUTPUT 1 2 21 6
c0 1 507 8.8e-13
c2 505 504 6e-14
c3 503 504 6e-14
d0 504 503 DSIM2
d1 505 504 DSIM2
d2 506 505 DSIM1
d3 503 501 DSIM1
e0 506 2 508 0 1
e1 6 501 502 0 1
e2 507 0 6 2 0.5
g0 0 505 VALUE = {LIMIT (-0.0042667*V(21,0),0.00032,-0.00032)}
g1 503 0 VALUE = {LIMIT (0.0042667*V(21,0),0.00032,-0.00032)}
g2 6 0 VALUE = {LIMIT (-0.0085333*V(21,0),0.00064,0)}
g3 0 2 VALUE = {LIMIT (0.0085333*V(21,0),0.00064,0)}
i4 0 508 dc 0.001
i5 0 502 dc 0.001
q0 504 505 2 2 NPN_OUT
q1 504 503 6 2 PNP_OUT
r0 1 507 50000
r1 504 1 10
r3 508 0 850 tc=-0.00302
r4 502 0 850 tc=-0.00302
.ENDS

*
* Models Used
*
.model DESD d cjo=5e-14 is=1e-17 rs=0.5 eg=1.12
.model DSIM1 d is=1e-12
.model DSIM2 d is=1e-14 eg=0.950
.model DSIM3 d is=1e-15
.model NPN_IN1 npn bf=140 cjc=1.20e-14 cje=2.78e-14 is=9.1e-18 rb=60 re=400 tf=4.7e-12
.model NPN_IN2 npn bf=1e6 cjc=1.20e-14 cje=2.78e-14 is=9.1e-18 rb=60 re=400 tf=4.7e-12
.model PNP_IN1 pnp bf=25 cjc=5.50e-14 cje=1.05e-13 is=3.5e-17 rb=75 re=600 tf=1.2e-12
.model NPN_OUT npn bf=75 cjc=1.60e-13 cjs=6.5e-14 is=1.0e-16 vaf=50
.model PNP_OUT pnp bf=60 cjc=1.50e-13 cjs=6.5e-14 is=6.4e-17 vaf=30