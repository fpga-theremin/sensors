/*********************************************/
/* SINE table of size 4096 and 13-bit values */
/* Latency: 4 CLK cycles                     */
/*********************************************/
module sin_cos_table_4096_13bit #(
    parameter DATA_WIDTH = 13,
    parameter ADDR_WIDTH = 12
)
(
    /* input clock                                           */
    input wire CLK,
    /* clock enable, 1 = enable pipeline, 0 = pause pipeline */
    input wire CE,
    /* reset signal, active 1                                */
    input wire RESET,
    
    /* sine table address to get value from                  */
    input wire [ADDR_WIDTH-1:0] PHASE,
    /* sin sample value from ROM, delayed by 4 clock cycles */
    output wire [DATA_WIDTH-1:0] SIN_VALUE,
    /* cos sample value from ROM, delayed by 4 clock cycles */
    output wire [DATA_WIDTH-1:0] COS_VALUE
    
);
    
    
    /* ROM size: we need to store only 1/4 of table entries, the rest may be obtained by mirroring and changing the sign */
    localparam MEMSIZE = 1 << (ADDR_WIDTH - 2);
    
    /* first quarter of table always has 0 in upper bit, so we can store only DATA_WIDTH-1 bits in the table */
    (* ram_style = "block" *)  
    reg [DATA_WIDTH-2:0] memory[0:MEMSIZE-1];
           
    /* store input phase value in register */
    reg [ADDR_WIDTH-1:0] phase_stage0;
    always @(posedge CLK)
        if (RESET)
            phase_stage0 <= 0;
        else if (CE)
            phase_stage0 <= PHASE;
     
    wire [1:0] sin_phase_top = phase_stage0[ADDR_WIDTH-1:ADDR_WIDTH-2];
    wire [1:0] cos_phase_top = phase_stage0[ADDR_WIDTH-1:ADDR_WIDTH-2] + 1;
     
    /* second half of table is the same as first, but negative */
    wire sin_need_sign_change = sin_phase_top[1];
    /* second and third quarters of table are mirrored by phase */
    wire sin_need_phase_inverse = sin_phase_top[0];
     
    /* second half of table is the same as first, but negative */
    wire cos_need_sign_change = cos_phase_top[1];
    /* second and third quarters of table are mirrored by phase */
    wire cos_need_phase_inverse = cos_phase_top[0];
     
    /* SIN: invert phase to have mirrored value */
    wire [ADDR_WIDTH-3:0] sin_table_entry_index = phase_stage0[ADDR_WIDTH-3:0] ^ { (ADDR_WIDTH-2) {sin_need_phase_inverse} };
    /* COS: invert phase to have mirrored value */
    wire [ADDR_WIDTH-3:0] cos_table_entry_index = phase_stage0[ADDR_WIDTH-3:0] ^ { (ADDR_WIDTH-2) {cos_need_phase_inverse} };
     
    /* propagate sign change flag to support negative values */
    reg sin_need_sign_change_stage1;
    reg cos_need_sign_change_stage1;
    reg sin_need_sign_change_stage2;
    reg cos_need_sign_change_stage2;
     
    always @(posedge CLK)
        if (CE) begin
            sin_need_sign_change_stage1 <= sin_need_sign_change;
            sin_need_sign_change_stage2 <= sin_need_sign_change_stage1;
            cos_need_sign_change_stage1 <= cos_need_sign_change;
            cos_need_sign_change_stage2 <= cos_need_sign_change_stage1;
        end
            
    /* SIN table: block RAM based ROM - first stage of pipeline */
    reg [DATA_WIDTH-2:0] sin_rddata_stage1;
    always @(posedge CLK)
        if (CE)
            sin_rddata_stage1 <= memory[sin_table_entry_index];
     
    /* COS table: block RAM based ROM - first stage of pipeline */
    reg [DATA_WIDTH-2:0] cos_rddata_stage1;
    always @(posedge CLK)
        if (CE)
            cos_rddata_stage1 <= memory[cos_table_entry_index];
     
    /* SIN table: block RAM based ROM - second stage of pipeline */
    reg [DATA_WIDTH-2:0] sin_rddata_stage2;
    always @(posedge CLK)
        if (CE)
            sin_rddata_stage2 <= sin_rddata_stage1;
     
    /* COS table: block RAM based ROM - second stage of pipeline */
    reg [DATA_WIDTH-2:0] cos_rddata_stage2;
    always @(posedge CLK)
        if (CE)
            cos_rddata_stage2 <= cos_rddata_stage1;
     
    /* SIN: this is output stage register, need sign bit as well */
    reg [DATA_WIDTH-1:0] sin_rddata_stage3;
    always @(posedge CLK)
        if (RESET)
            sin_rddata_stage3 <= 0; 
        else if (CE)
            sin_rddata_stage3 <= sin_need_sign_change_stage2 ? -{1'b0, sin_rddata_stage2} : {1'b0, sin_rddata_stage2}; 
     
    /* COS: this is output stage register, need sign bit as well */
    reg [DATA_WIDTH-1:0] cos_rddata_stage3;
    always @(posedge CLK)
        if (RESET)
            cos_rddata_stage3 <= 0; 
        else if (CE)
            cos_rddata_stage3 <= cos_need_sign_change_stage2 ? -{1'b0, cos_rddata_stage2} : {1'b0, cos_rddata_stage2}; 
     
    /* propagate value to output */
    assign SIN_VALUE = sin_rddata_stage3;
    assign COS_VALUE = cos_rddata_stage3;
    
    

    /* Initialization of ROM content with first quarter of SINE function */
    initial begin
        memory[0] = 3;
        memory[1] = 9;
        memory[2] = 16;
        memory[3] = 22;
        memory[4] = 28;
        memory[5] = 35;
        memory[6] = 41;
        memory[7] = 47;
        memory[8] = 53;
        memory[9] = 60;
        memory[10] = 66;
        memory[11] = 72;
        memory[12] = 79;
        memory[13] = 85;
        memory[14] = 91;
        memory[15] = 97;
        memory[16] = 104;
        memory[17] = 110;
        memory[18] = 116;
        memory[19] = 122;
        memory[20] = 129;
        memory[21] = 135;
        memory[22] = 141;
        memory[23] = 148;
        memory[24] = 154;
        memory[25] = 160;
        memory[26] = 166;
        memory[27] = 173;
        memory[28] = 179;
        memory[29] = 185;
        memory[30] = 192;
        memory[31] = 198;
        memory[32] = 204;
        memory[33] = 210;
        memory[34] = 217;
        memory[35] = 223;
        memory[36] = 229;
        memory[37] = 235;
        memory[38] = 242;
        memory[39] = 248;
        memory[40] = 254;
        memory[41] = 261;
        memory[42] = 267;
        memory[43] = 273;
        memory[44] = 279;
        memory[45] = 286;
        memory[46] = 292;
        memory[47] = 298;
        memory[48] = 304;
        memory[49] = 311;
        memory[50] = 317;
        memory[51] = 323;
        memory[52] = 329;
        memory[53] = 336;
        memory[54] = 342;
        memory[55] = 348;
        memory[56] = 354;
        memory[57] = 361;
        memory[58] = 367;
        memory[59] = 373;
        memory[60] = 379;
        memory[61] = 386;
        memory[62] = 392;
        memory[63] = 398;
        memory[64] = 405;
        memory[65] = 411;
        memory[66] = 417;
        memory[67] = 423;
        memory[68] = 430;
        memory[69] = 436;
        memory[70] = 442;
        memory[71] = 448;
        memory[72] = 454;
        memory[73] = 461;
        memory[74] = 467;
        memory[75] = 473;
        memory[76] = 479;
        memory[77] = 486;
        memory[78] = 492;
        memory[79] = 498;
        memory[80] = 504;
        memory[81] = 511;
        memory[82] = 517;
        memory[83] = 523;
        memory[84] = 529;
        memory[85] = 536;
        memory[86] = 542;
        memory[87] = 548;
        memory[88] = 554;
        memory[89] = 560;
        memory[90] = 567;
        memory[91] = 573;
        memory[92] = 579;
        memory[93] = 585;
        memory[94] = 592;
        memory[95] = 598;
        memory[96] = 604;
        memory[97] = 610;
        memory[98] = 616;
        memory[99] = 623;
        memory[100] = 629;
        memory[101] = 635;
        memory[102] = 641;
        memory[103] = 647;
        memory[104] = 654;
        memory[105] = 660;
        memory[106] = 666;
        memory[107] = 672;
        memory[108] = 678;
        memory[109] = 685;
        memory[110] = 691;
        memory[111] = 697;
        memory[112] = 703;
        memory[113] = 709;
        memory[114] = 716;
        memory[115] = 722;
        memory[116] = 728;
        memory[117] = 734;
        memory[118] = 740;
        memory[119] = 746;
        memory[120] = 753;
        memory[121] = 759;
        memory[122] = 765;
        memory[123] = 771;
        memory[124] = 777;
        memory[125] = 783;
        memory[126] = 790;
        memory[127] = 796;
        memory[128] = 802;
        memory[129] = 808;
        memory[130] = 814;
        memory[131] = 820;
        memory[132] = 827;
        memory[133] = 833;
        memory[134] = 839;
        memory[135] = 845;
        memory[136] = 851;
        memory[137] = 857;
        memory[138] = 863;
        memory[139] = 870;
        memory[140] = 876;
        memory[141] = 882;
        memory[142] = 888;
        memory[143] = 894;
        memory[144] = 900;
        memory[145] = 906;
        memory[146] = 913;
        memory[147] = 919;
        memory[148] = 925;
        memory[149] = 931;
        memory[150] = 937;
        memory[151] = 943;
        memory[152] = 949;
        memory[153] = 955;
        memory[154] = 961;
        memory[155] = 968;
        memory[156] = 974;
        memory[157] = 980;
        memory[158] = 986;
        memory[159] = 992;
        memory[160] = 998;
        memory[161] = 1004;
        memory[162] = 1010;
        memory[163] = 1016;
        memory[164] = 1022;
        memory[165] = 1028;
        memory[166] = 1035;
        memory[167] = 1041;
        memory[168] = 1047;
        memory[169] = 1053;
        memory[170] = 1059;
        memory[171] = 1065;
        memory[172] = 1071;
        memory[173] = 1077;
        memory[174] = 1083;
        memory[175] = 1089;
        memory[176] = 1095;
        memory[177] = 1101;
        memory[178] = 1107;
        memory[179] = 1113;
        memory[180] = 1119;
        memory[181] = 1125;
        memory[182] = 1131;
        memory[183] = 1138;
        memory[184] = 1144;
        memory[185] = 1150;
        memory[186] = 1156;
        memory[187] = 1162;
        memory[188] = 1168;
        memory[189] = 1174;
        memory[190] = 1180;
        memory[191] = 1186;
        memory[192] = 1192;
        memory[193] = 1198;
        memory[194] = 1204;
        memory[195] = 1210;
        memory[196] = 1216;
        memory[197] = 1222;
        memory[198] = 1228;
        memory[199] = 1234;
        memory[200] = 1240;
        memory[201] = 1246;
        memory[202] = 1252;
        memory[203] = 1258;
        memory[204] = 1264;
        memory[205] = 1270;
        memory[206] = 1276;
        memory[207] = 1282;
        memory[208] = 1288;
        memory[209] = 1293;
        memory[210] = 1299;
        memory[211] = 1305;
        memory[212] = 1311;
        memory[213] = 1317;
        memory[214] = 1323;
        memory[215] = 1329;
        memory[216] = 1335;
        memory[217] = 1341;
        memory[218] = 1347;
        memory[219] = 1353;
        memory[220] = 1359;
        memory[221] = 1365;
        memory[222] = 1371;
        memory[223] = 1377;
        memory[224] = 1383;
        memory[225] = 1388;
        memory[226] = 1394;
        memory[227] = 1400;
        memory[228] = 1406;
        memory[229] = 1412;
        memory[230] = 1418;
        memory[231] = 1424;
        memory[232] = 1430;
        memory[233] = 1436;
        memory[234] = 1441;
        memory[235] = 1447;
        memory[236] = 1453;
        memory[237] = 1459;
        memory[238] = 1465;
        memory[239] = 1471;
        memory[240] = 1477;
        memory[241] = 1483;
        memory[242] = 1488;
        memory[243] = 1494;
        memory[244] = 1500;
        memory[245] = 1506;
        memory[246] = 1512;
        memory[247] = 1518;
        memory[248] = 1523;
        memory[249] = 1529;
        memory[250] = 1535;
        memory[251] = 1541;
        memory[252] = 1547;
        memory[253] = 1553;
        memory[254] = 1558;
        memory[255] = 1564;
        memory[256] = 1570;
        memory[257] = 1576;
        memory[258] = 1582;
        memory[259] = 1587;
        memory[260] = 1593;
        memory[261] = 1599;
        memory[262] = 1605;
        memory[263] = 1611;
        memory[264] = 1616;
        memory[265] = 1622;
        memory[266] = 1628;
        memory[267] = 1634;
        memory[268] = 1639;
        memory[269] = 1645;
        memory[270] = 1651;
        memory[271] = 1657;
        memory[272] = 1662;
        memory[273] = 1668;
        memory[274] = 1674;
        memory[275] = 1680;
        memory[276] = 1685;
        memory[277] = 1691;
        memory[278] = 1697;
        memory[279] = 1702;
        memory[280] = 1708;
        memory[281] = 1714;
        memory[282] = 1720;
        memory[283] = 1725;
        memory[284] = 1731;
        memory[285] = 1737;
        memory[286] = 1742;
        memory[287] = 1748;
        memory[288] = 1754;
        memory[289] = 1759;
        memory[290] = 1765;
        memory[291] = 1771;
        memory[292] = 1776;
        memory[293] = 1782;
        memory[294] = 1788;
        memory[295] = 1793;
        memory[296] = 1799;
        memory[297] = 1805;
        memory[298] = 1810;
        memory[299] = 1816;
        memory[300] = 1821;
        memory[301] = 1827;
        memory[302] = 1833;
        memory[303] = 1838;
        memory[304] = 1844;
        memory[305] = 1850;
        memory[306] = 1855;
        memory[307] = 1861;
        memory[308] = 1866;
        memory[309] = 1872;
        memory[310] = 1878;
        memory[311] = 1883;
        memory[312] = 1889;
        memory[313] = 1894;
        memory[314] = 1900;
        memory[315] = 1905;
        memory[316] = 1911;
        memory[317] = 1917;
        memory[318] = 1922;
        memory[319] = 1928;
        memory[320] = 1933;
        memory[321] = 1939;
        memory[322] = 1944;
        memory[323] = 1950;
        memory[324] = 1955;
        memory[325] = 1961;
        memory[326] = 1966;
        memory[327] = 1972;
        memory[328] = 1977;
        memory[329] = 1983;
        memory[330] = 1988;
        memory[331] = 1994;
        memory[332] = 1999;
        memory[333] = 2005;
        memory[334] = 2010;
        memory[335] = 2016;
        memory[336] = 2021;
        memory[337] = 2027;
        memory[338] = 2032;
        memory[339] = 2038;
        memory[340] = 2043;
        memory[341] = 2048;
        memory[342] = 2054;
        memory[343] = 2059;
        memory[344] = 2065;
        memory[345] = 2070;
        memory[346] = 2076;
        memory[347] = 2081;
        memory[348] = 2086;
        memory[349] = 2092;
        memory[350] = 2097;
        memory[351] = 2103;
        memory[352] = 2108;
        memory[353] = 2113;
        memory[354] = 2119;
        memory[355] = 2124;
        memory[356] = 2129;
        memory[357] = 2135;
        memory[358] = 2140;
        memory[359] = 2146;
        memory[360] = 2151;
        memory[361] = 2156;
        memory[362] = 2162;
        memory[363] = 2167;
        memory[364] = 2172;
        memory[365] = 2178;
        memory[366] = 2183;
        memory[367] = 2188;
        memory[368] = 2193;
        memory[369] = 2199;
        memory[370] = 2204;
        memory[371] = 2209;
        memory[372] = 2215;
        memory[373] = 2220;
        memory[374] = 2225;
        memory[375] = 2230;
        memory[376] = 2236;
        memory[377] = 2241;
        memory[378] = 2246;
        memory[379] = 2252;
        memory[380] = 2257;
        memory[381] = 2262;
        memory[382] = 2267;
        memory[383] = 2272;
        memory[384] = 2278;
        memory[385] = 2283;
        memory[386] = 2288;
        memory[387] = 2293;
        memory[388] = 2299;
        memory[389] = 2304;
        memory[390] = 2309;
        memory[391] = 2314;
        memory[392] = 2319;
        memory[393] = 2324;
        memory[394] = 2330;
        memory[395] = 2335;
        memory[396] = 2340;
        memory[397] = 2345;
        memory[398] = 2350;
        memory[399] = 2355;
        memory[400] = 2361;
        memory[401] = 2366;
        memory[402] = 2371;
        memory[403] = 2376;
        memory[404] = 2381;
        memory[405] = 2386;
        memory[406] = 2391;
        memory[407] = 2396;
        memory[408] = 2401;
        memory[409] = 2406;
        memory[410] = 2412;
        memory[411] = 2417;
        memory[412] = 2422;
        memory[413] = 2427;
        memory[414] = 2432;
        memory[415] = 2437;
        memory[416] = 2442;
        memory[417] = 2447;
        memory[418] = 2452;
        memory[419] = 2457;
        memory[420] = 2462;
        memory[421] = 2467;
        memory[422] = 2472;
        memory[423] = 2477;
        memory[424] = 2482;
        memory[425] = 2487;
        memory[426] = 2492;
        memory[427] = 2497;
        memory[428] = 2502;
        memory[429] = 2507;
        memory[430] = 2512;
        memory[431] = 2517;
        memory[432] = 2522;
        memory[433] = 2527;
        memory[434] = 2532;
        memory[435] = 2537;
        memory[436] = 2542;
        memory[437] = 2547;
        memory[438] = 2551;
        memory[439] = 2556;
        memory[440] = 2561;
        memory[441] = 2566;
        memory[442] = 2571;
        memory[443] = 2576;
        memory[444] = 2581;
        memory[445] = 2586;
        memory[446] = 2591;
        memory[447] = 2595;
        memory[448] = 2600;
        memory[449] = 2605;
        memory[450] = 2610;
        memory[451] = 2615;
        memory[452] = 2620;
        memory[453] = 2624;
        memory[454] = 2629;
        memory[455] = 2634;
        memory[456] = 2639;
        memory[457] = 2644;
        memory[458] = 2648;
        memory[459] = 2653;
        memory[460] = 2658;
        memory[461] = 2663;
        memory[462] = 2668;
        memory[463] = 2672;
        memory[464] = 2677;
        memory[465] = 2682;
        memory[466] = 2687;
        memory[467] = 2691;
        memory[468] = 2696;
        memory[469] = 2701;
        memory[470] = 2706;
        memory[471] = 2710;
        memory[472] = 2715;
        memory[473] = 2720;
        memory[474] = 2724;
        memory[475] = 2729;
        memory[476] = 2734;
        memory[477] = 2738;
        memory[478] = 2743;
        memory[479] = 2748;
        memory[480] = 2752;
        memory[481] = 2757;
        memory[482] = 2762;
        memory[483] = 2766;
        memory[484] = 2771;
        memory[485] = 2776;
        memory[486] = 2780;
        memory[487] = 2785;
        memory[488] = 2789;
        memory[489] = 2794;
        memory[490] = 2799;
        memory[491] = 2803;
        memory[492] = 2808;
        memory[493] = 2812;
        memory[494] = 2817;
        memory[495] = 2821;
        memory[496] = 2826;
        memory[497] = 2830;
        memory[498] = 2835;
        memory[499] = 2840;
        memory[500] = 2844;
        memory[501] = 2849;
        memory[502] = 2853;
        memory[503] = 2858;
        memory[504] = 2862;
        memory[505] = 2867;
        memory[506] = 2871;
        memory[507] = 2876;
        memory[508] = 2880;
        memory[509] = 2884;
        memory[510] = 2889;
        memory[511] = 2893;
        memory[512] = 2898;
        memory[513] = 2902;
        memory[514] = 2907;
        memory[515] = 2911;
        memory[516] = 2916;
        memory[517] = 2920;
        memory[518] = 2924;
        memory[519] = 2929;
        memory[520] = 2933;
        memory[521] = 2937;
        memory[522] = 2942;
        memory[523] = 2946;
        memory[524] = 2951;
        memory[525] = 2955;
        memory[526] = 2959;
        memory[527] = 2964;
        memory[528] = 2968;
        memory[529] = 2972;
        memory[530] = 2977;
        memory[531] = 2981;
        memory[532] = 2985;
        memory[533] = 2990;
        memory[534] = 2994;
        memory[535] = 2998;
        memory[536] = 3002;
        memory[537] = 3007;
        memory[538] = 3011;
        memory[539] = 3015;
        memory[540] = 3019;
        memory[541] = 3024;
        memory[542] = 3028;
        memory[543] = 3032;
        memory[544] = 3036;
        memory[545] = 3041;
        memory[546] = 3045;
        memory[547] = 3049;
        memory[548] = 3053;
        memory[549] = 3057;
        memory[550] = 3061;
        memory[551] = 3066;
        memory[552] = 3070;
        memory[553] = 3074;
        memory[554] = 3078;
        memory[555] = 3082;
        memory[556] = 3086;
        memory[557] = 3090;
        memory[558] = 3095;
        memory[559] = 3099;
        memory[560] = 3103;
        memory[561] = 3107;
        memory[562] = 3111;
        memory[563] = 3115;
        memory[564] = 3119;
        memory[565] = 3123;
        memory[566] = 3127;
        memory[567] = 3131;
        memory[568] = 3135;
        memory[569] = 3139;
        memory[570] = 3143;
        memory[571] = 3147;
        memory[572] = 3151;
        memory[573] = 3155;
        memory[574] = 3159;
        memory[575] = 3163;
        memory[576] = 3167;
        memory[577] = 3171;
        memory[578] = 3175;
        memory[579] = 3179;
        memory[580] = 3183;
        memory[581] = 3187;
        memory[582] = 3191;
        memory[583] = 3195;
        memory[584] = 3199;
        memory[585] = 3203;
        memory[586] = 3207;
        memory[587] = 3211;
        memory[588] = 3215;
        memory[589] = 3219;
        memory[590] = 3222;
        memory[591] = 3226;
        memory[592] = 3230;
        memory[593] = 3234;
        memory[594] = 3238;
        memory[595] = 3242;
        memory[596] = 3246;
        memory[597] = 3249;
        memory[598] = 3253;
        memory[599] = 3257;
        memory[600] = 3261;
        memory[601] = 3265;
        memory[602] = 3268;
        memory[603] = 3272;
        memory[604] = 3276;
        memory[605] = 3280;
        memory[606] = 3284;
        memory[607] = 3287;
        memory[608] = 3291;
        memory[609] = 3295;
        memory[610] = 3298;
        memory[611] = 3302;
        memory[612] = 3306;
        memory[613] = 3310;
        memory[614] = 3313;
        memory[615] = 3317;
        memory[616] = 3321;
        memory[617] = 3324;
        memory[618] = 3328;
        memory[619] = 3332;
        memory[620] = 3335;
        memory[621] = 3339;
        memory[622] = 3343;
        memory[623] = 3346;
        memory[624] = 3350;
        memory[625] = 3353;
        memory[626] = 3357;
        memory[627] = 3361;
        memory[628] = 3364;
        memory[629] = 3368;
        memory[630] = 3371;
        memory[631] = 3375;
        memory[632] = 3378;
        memory[633] = 3382;
        memory[634] = 3386;
        memory[635] = 3389;
        memory[636] = 3393;
        memory[637] = 3396;
        memory[638] = 3400;
        memory[639] = 3403;
        memory[640] = 3407;
        memory[641] = 3410;
        memory[642] = 3414;
        memory[643] = 3417;
        memory[644] = 3420;
        memory[645] = 3424;
        memory[646] = 3427;
        memory[647] = 3431;
        memory[648] = 3434;
        memory[649] = 3438;
        memory[650] = 3441;
        memory[651] = 3444;
        memory[652] = 3448;
        memory[653] = 3451;
        memory[654] = 3455;
        memory[655] = 3458;
        memory[656] = 3461;
        memory[657] = 3465;
        memory[658] = 3468;
        memory[659] = 3471;
        memory[660] = 3475;
        memory[661] = 3478;
        memory[662] = 3481;
        memory[663] = 3485;
        memory[664] = 3488;
        memory[665] = 3491;
        memory[666] = 3495;
        memory[667] = 3498;
        memory[668] = 3501;
        memory[669] = 3504;
        memory[670] = 3508;
        memory[671] = 3511;
        memory[672] = 3514;
        memory[673] = 3517;
        memory[674] = 3520;
        memory[675] = 3524;
        memory[676] = 3527;
        memory[677] = 3530;
        memory[678] = 3533;
        memory[679] = 3536;
        memory[680] = 3540;
        memory[681] = 3543;
        memory[682] = 3546;
        memory[683] = 3549;
        memory[684] = 3552;
        memory[685] = 3555;
        memory[686] = 3558;
        memory[687] = 3561;
        memory[688] = 3565;
        memory[689] = 3568;
        memory[690] = 3571;
        memory[691] = 3574;
        memory[692] = 3577;
        memory[693] = 3580;
        memory[694] = 3583;
        memory[695] = 3586;
        memory[696] = 3589;
        memory[697] = 3592;
        memory[698] = 3595;
        memory[699] = 3598;
        memory[700] = 3601;
        memory[701] = 3604;
        memory[702] = 3607;
        memory[703] = 3610;
        memory[704] = 3613;
        memory[705] = 3616;
        memory[706] = 3619;
        memory[707] = 3622;
        memory[708] = 3625;
        memory[709] = 3628;
        memory[710] = 3631;
        memory[711] = 3633;
        memory[712] = 3636;
        memory[713] = 3639;
        memory[714] = 3642;
        memory[715] = 3645;
        memory[716] = 3648;
        memory[717] = 3651;
        memory[718] = 3654;
        memory[719] = 3656;
        memory[720] = 3659;
        memory[721] = 3662;
        memory[722] = 3665;
        memory[723] = 3668;
        memory[724] = 3670;
        memory[725] = 3673;
        memory[726] = 3676;
        memory[727] = 3679;
        memory[728] = 3681;
        memory[729] = 3684;
        memory[730] = 3687;
        memory[731] = 3690;
        memory[732] = 3692;
        memory[733] = 3695;
        memory[734] = 3698;
        memory[735] = 3700;
        memory[736] = 3703;
        memory[737] = 3706;
        memory[738] = 3709;
        memory[739] = 3711;
        memory[740] = 3714;
        memory[741] = 3716;
        memory[742] = 3719;
        memory[743] = 3722;
        memory[744] = 3724;
        memory[745] = 3727;
        memory[746] = 3730;
        memory[747] = 3732;
        memory[748] = 3735;
        memory[749] = 3737;
        memory[750] = 3740;
        memory[751] = 3742;
        memory[752] = 3745;
        memory[753] = 3747;
        memory[754] = 3750;
        memory[755] = 3753;
        memory[756] = 3755;
        memory[757] = 3758;
        memory[758] = 3760;
        memory[759] = 3763;
        memory[760] = 3765;
        memory[761] = 3767;
        memory[762] = 3770;
        memory[763] = 3772;
        memory[764] = 3775;
        memory[765] = 3777;
        memory[766] = 3780;
        memory[767] = 3782;
        memory[768] = 3784;
        memory[769] = 3787;
        memory[770] = 3789;
        memory[771] = 3792;
        memory[772] = 3794;
        memory[773] = 3796;
        memory[774] = 3799;
        memory[775] = 3801;
        memory[776] = 3803;
        memory[777] = 3806;
        memory[778] = 3808;
        memory[779] = 3810;
        memory[780] = 3813;
        memory[781] = 3815;
        memory[782] = 3817;
        memory[783] = 3819;
        memory[784] = 3822;
        memory[785] = 3824;
        memory[786] = 3826;
        memory[787] = 3828;
        memory[788] = 3831;
        memory[789] = 3833;
        memory[790] = 3835;
        memory[791] = 3837;
        memory[792] = 3839;
        memory[793] = 3842;
        memory[794] = 3844;
        memory[795] = 3846;
        memory[796] = 3848;
        memory[797] = 3850;
        memory[798] = 3852;
        memory[799] = 3855;
        memory[800] = 3857;
        memory[801] = 3859;
        memory[802] = 3861;
        memory[803] = 3863;
        memory[804] = 3865;
        memory[805] = 3867;
        memory[806] = 3869;
        memory[807] = 3871;
        memory[808] = 3873;
        memory[809] = 3875;
        memory[810] = 3877;
        memory[811] = 3879;
        memory[812] = 3881;
        memory[813] = 3883;
        memory[814] = 3885;
        memory[815] = 3887;
        memory[816] = 3889;
        memory[817] = 3891;
        memory[818] = 3893;
        memory[819] = 3895;
        memory[820] = 3897;
        memory[821] = 3899;
        memory[822] = 3901;
        memory[823] = 3903;
        memory[824] = 3905;
        memory[825] = 3907;
        memory[826] = 3909;
        memory[827] = 3910;
        memory[828] = 3912;
        memory[829] = 3914;
        memory[830] = 3916;
        memory[831] = 3918;
        memory[832] = 3920;
        memory[833] = 3921;
        memory[834] = 3923;
        memory[835] = 3925;
        memory[836] = 3927;
        memory[837] = 3929;
        memory[838] = 3930;
        memory[839] = 3932;
        memory[840] = 3934;
        memory[841] = 3936;
        memory[842] = 3937;
        memory[843] = 3939;
        memory[844] = 3941;
        memory[845] = 3942;
        memory[846] = 3944;
        memory[847] = 3946;
        memory[848] = 3947;
        memory[849] = 3949;
        memory[850] = 3951;
        memory[851] = 3952;
        memory[852] = 3954;
        memory[853] = 3956;
        memory[854] = 3957;
        memory[855] = 3959;
        memory[856] = 3961;
        memory[857] = 3962;
        memory[858] = 3964;
        memory[859] = 3965;
        memory[860] = 3967;
        memory[861] = 3968;
        memory[862] = 3970;
        memory[863] = 3972;
        memory[864] = 3973;
        memory[865] = 3975;
        memory[866] = 3976;
        memory[867] = 3978;
        memory[868] = 3979;
        memory[869] = 3981;
        memory[870] = 3982;
        memory[871] = 3983;
        memory[872] = 3985;
        memory[873] = 3986;
        memory[874] = 3988;
        memory[875] = 3989;
        memory[876] = 3991;
        memory[877] = 3992;
        memory[878] = 3993;
        memory[879] = 3995;
        memory[880] = 3996;
        memory[881] = 3998;
        memory[882] = 3999;
        memory[883] = 4000;
        memory[884] = 4002;
        memory[885] = 4003;
        memory[886] = 4004;
        memory[887] = 4006;
        memory[888] = 4007;
        memory[889] = 4008;
        memory[890] = 4009;
        memory[891] = 4011;
        memory[892] = 4012;
        memory[893] = 4013;
        memory[894] = 4014;
        memory[895] = 4016;
        memory[896] = 4017;
        memory[897] = 4018;
        memory[898] = 4019;
        memory[899] = 4021;
        memory[900] = 4022;
        memory[901] = 4023;
        memory[902] = 4024;
        memory[903] = 4025;
        memory[904] = 4026;
        memory[905] = 4028;
        memory[906] = 4029;
        memory[907] = 4030;
        memory[908] = 4031;
        memory[909] = 4032;
        memory[910] = 4033;
        memory[911] = 4034;
        memory[912] = 4035;
        memory[913] = 4036;
        memory[914] = 4037;
        memory[915] = 4038;
        memory[916] = 4039;
        memory[917] = 4040;
        memory[918] = 4041;
        memory[919] = 4042;
        memory[920] = 4043;
        memory[921] = 4044;
        memory[922] = 4045;
        memory[923] = 4046;
        memory[924] = 4047;
        memory[925] = 4048;
        memory[926] = 4049;
        memory[927] = 4050;
        memory[928] = 4051;
        memory[929] = 4052;
        memory[930] = 4053;
        memory[931] = 4054;
        memory[932] = 4055;
        memory[933] = 4056;
        memory[934] = 4056;
        memory[935] = 4057;
        memory[936] = 4058;
        memory[937] = 4059;
        memory[938] = 4060;
        memory[939] = 4061;
        memory[940] = 4061;
        memory[941] = 4062;
        memory[942] = 4063;
        memory[943] = 4064;
        memory[944] = 4065;
        memory[945] = 4065;
        memory[946] = 4066;
        memory[947] = 4067;
        memory[948] = 4068;
        memory[949] = 4068;
        memory[950] = 4069;
        memory[951] = 4070;
        memory[952] = 4070;
        memory[953] = 4071;
        memory[954] = 4072;
        memory[955] = 4072;
        memory[956] = 4073;
        memory[957] = 4074;
        memory[958] = 4074;
        memory[959] = 4075;
        memory[960] = 4076;
        memory[961] = 4076;
        memory[962] = 4077;
        memory[963] = 4077;
        memory[964] = 4078;
        memory[965] = 4079;
        memory[966] = 4079;
        memory[967] = 4080;
        memory[968] = 4080;
        memory[969] = 4081;
        memory[970] = 4081;
        memory[971] = 4082;
        memory[972] = 4082;
        memory[973] = 4083;
        memory[974] = 4083;
        memory[975] = 4084;
        memory[976] = 4084;
        memory[977] = 4085;
        memory[978] = 4085;
        memory[979] = 4085;
        memory[980] = 4086;
        memory[981] = 4086;
        memory[982] = 4087;
        memory[983] = 4087;
        memory[984] = 4087;
        memory[985] = 4088;
        memory[986] = 4088;
        memory[987] = 4089;
        memory[988] = 4089;
        memory[989] = 4089;
        memory[990] = 4090;
        memory[991] = 4090;
        memory[992] = 4090;
        memory[993] = 4091;
        memory[994] = 4091;
        memory[995] = 4091;
        memory[996] = 4091;
        memory[997] = 4092;
        memory[998] = 4092;
        memory[999] = 4092;
        memory[1000] = 4092;
        memory[1001] = 4093;
        memory[1002] = 4093;
        memory[1003] = 4093;
        memory[1004] = 4093;
        memory[1005] = 4093;
        memory[1006] = 4094;
        memory[1007] = 4094;
        memory[1008] = 4094;
        memory[1009] = 4094;
        memory[1010] = 4094;
        memory[1011] = 4094;
        memory[1012] = 4094;
        memory[1013] = 4094;
        memory[1014] = 4095;
        memory[1015] = 4095;
        memory[1016] = 4095;
        memory[1017] = 4095;
        memory[1018] = 4095;
        memory[1019] = 4095;
        memory[1020] = 4095;
        memory[1021] = 4095;
        memory[1022] = 4095;
        memory[1023] = 4095;
    end

endmodule
